Borehole ID|CampCentury
Place name|Camp Century
Geographic location|Northwest Greenland
Site type|Ice sheet
Data Source|Graphic in science source
Data DOI|
Science Source|Gundestrup, N. S., Dahl-Jensen, D., Hansen, B. L., & Kelty, J. (1993). Bore-hole survey at Camp Century, 1989. Cold regions science and technology, 21(2), 187-193.
Science DOI|10.1016/0165-232X(93)90006-T
Date|1966
Longitude [°E]|-61.1097
Latitude [°N]|77.1797
Location Source|Colgan, 2021
Depth of top measurement [m]|100.0
Depth of bottom measurement [m]|1387
Ice thickness [m]|1387
Coverage [% of thickness]|93
Ice thickness source|Weertman, 1968
Note|Data from Gundestrup (1993) seems higher fidelity than Weertman (1968). See https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/issues/38
