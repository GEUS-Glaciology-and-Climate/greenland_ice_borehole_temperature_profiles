Name|agassiz79a
Alternate name|Agassiz ice cap 1979A borehole 
Data source|WIC Email 
Drill year(s)|nan 
Data year(s)|1979 
Longitude [°E]|-73.1 
Latitude [°N]|80.7 
Approximate location name|Agassiz Ice Cap 
Location source|See data source 
Ice thickness [m]|141.9 
Ice thickness year|nan 
Ice thickness source|See data source 
Surface velocity [m yr^-1]|nan 
Surface velocity year|nan 
Surface velocity source|nan 
Measured from: Top, Bottom, Relative|T 
Depth of top measurement [m]|12.0 
Depth of bottom measurement [m]|142.0 
Coverage [% of thickness]|92 
