Borehole ID|Isunnguata_27km-11B
Place Name|Isunnguata Sermia
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|T. Meierbachtol email
Data DOI|
Science Reference|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A943
Date|2011
Longitude [°E]|-49.71913
Latitude [°N]|67.19527
Location source|T. Meierbachtol email
Depth of top measurement [m]|27.0
Depth of bottom measurement [m]|460.0
Ice thickness [m]|466
Coverage [% of thickness]|93
Ice thickness source|T. Meierbachtol email
Measured from: Top, Bottom, Relative|T
General_Note|See data in M1-10 folder
Temperature_note|
Thickness_note|
Location_note|Harrington 2015 name: S3-B
