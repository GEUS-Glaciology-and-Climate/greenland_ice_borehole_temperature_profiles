Borehole ID|Meighen67
Place Name|Meighen Ice Cap
Geographic Location|Canadian Arctic North
Ice Type|Ice sheet
Data Reference|Paterson, W. S. B.: A temperature profile through the Meighen ice cap, Arctic Canada , International Association of Scientific Hydrology 79, 440–449, 1968 
Data DOI|
Science Reference|Paterson, W. S. B.: A temperature profile through the Meighen ice cap, Arctic Canada , International Association of Scientific Hydrology 79, 440–449, 1968 
Science DOI|
Date|1965
Longitude [°E]|-99.1
Latitude [°N]|79.9
Location source|See data source
Depth of top measurement [m]|1.0
Depth of bottom measurement [m]|121
Ice thickness [m]|121.2
Coverage [% of thickness]|99
Ice thickness source|See data source
General_Note|
Temperature_note|
Thickness_note|
Location_note|Location from Geothermal Database
