Borehole ID|CampVI
Place Name|Camp VI
Geographic Location|Central West Greenland
Ice Type|Sheet -Main
Data Reference|Digitization from published graphic
Data DOI|
Science Reference|
Science DOI|
Date|1950
Longitude [°E]|-48.2625
Latitude [°N]|69.6981
Location source|Heuberger1954
Depth of top measurement [m]|4.0
Depth of bottom measurement [m]|125.0
Ice thickness [m]|1389.0
Coverage [% of thickness]|9
Ice thickness source|BedMachine_V3
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
