Borehole ID|HansTausen_Hare
Place name|Hans Tausen Hare
Geographic location|North Greenland
Ice type|Ice cap
Data Source|Zekollari email
Data DOI|
Science Source|Thomsen, H., Reeh, N., Olesen, O., & Jonsson, P. (1996). Glacier and climate research on Hans Tausen Iskappe, North Greenland – 1995 glacier basin activities and preliminary results. Bulletin Grønlands Geologiske Undersøgelse, 172, 78–84. https://doi.org/10.34194/bullggu.v172.6749
Science DOI|10.34194/bullggu.v172.6749
Date|1995
Longitude [°E]|-36.67
Latitude [°N]|82.84
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|9.0
Depth of bottom measurement [m]|288
Ice thickness [m]|289
Coverage [% of thickness]|97
Ice thickness source|See data source
Note|Drill date: 10.34194/bullggu.v172.6749 
