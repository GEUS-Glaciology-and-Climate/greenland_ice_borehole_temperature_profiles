Borehole ID|FOXX1
Place name|Sermeq Avannerleq
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Ryser, C., Lüthi, M. P., Andrews, L. C., Hoffman, M. J., Catania, G. A., Hawley, R. L., ... & Kristensen, S. S. (2014). Sustained high basal motion of the Greenland ice sheet revealed by borehole deformation. Journal of Glaciology, 60(222), 647-660.
Data DOI|10.3189/2014JoG13J196
Science Source|Ryser, C., Lüthi, M. P., Andrews, L. C., Hoffman, M. J., Catania, G. A., Hawley, R. L., ... & Kristensen, S. S. (2014). Sustained high basal motion of the Greenland ice sheet revealed by borehole deformation. Journal of Glaciology, 60(222), 647-660.
Science DOI|10.3189/2014JoG13J196
Date|2012
Longitude [°E]|-49.8851
Latitude [°N]|69.4459
Location Source|10.3189/2014JoG13J196
Depth of top measurement [m]|411.0
Depth of bottom measurement [m]|606
Ice thickness [m]|624
Coverage [% of thickness]|31
Ice thickness source|Ryser, 2014 (Table 2)
Note|Date: Data was collected in 2011 and 2012 and the data extracted from the cooling curves
