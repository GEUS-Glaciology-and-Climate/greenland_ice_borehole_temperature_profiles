Borehole ID|GULL
Place name|Sermeq Avannerleq
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Graphic in science source
Data DOI|
Science Source|Lüthi, M., C. Ryser, L. Andrews et al. 2015. Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming. The Cryosphere. 9: 245-253. 
Science DOI|10.5194/tc-9-245-2015
Date|2012
Longitude [°E]|-49.7142
Latitude [°N]|69.4526
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|4.0
Depth of bottom measurement [m]|704
Ice thickness [m]|703
Coverage [% of thickness]|100
Ice thickness source|See data source
Note|Location from Geothermal Database; Date: Data was collected in 2011 and 2012 and the data extracted from the cooling curves
