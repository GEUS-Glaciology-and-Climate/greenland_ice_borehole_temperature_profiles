Borehole ID|td42
Descriptive Name|
Area|Paakitsoq
Data reference|Unknown PDF: See td1
Data DOI|
Science reference|
Science DOI|
Date|1991-08-28
Longitude [°E]|-49.683
Latitude [°N]|69.533
Location source|Unknown PDF: See td1
Depth of top measurement [m]|3.0
Depth of bottom measurement [m]|493.0
Ice thickness [m]|>600
Coverage [% of thickness]|#VALUE!
Ice thickness source|Unknown PDF: See td1
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
