Borehole ID|doyle_2018
Descriptive Name|
Area|Store Glacier
Data reference|Doyle, Samuel; Hubbard, Bryn; Christoffersen, Poul; Young, Tun Jan; Hofstede, Coen; Bougamont, Marion; et al. (2018): SAFIRE borehole, AWS and GPS datasets. figshare. Dataset. https://doi.org/10.6084/m9.figshare.5745294.v1 
Data DOI|10.6084/m9.figshare.5745294.v1
Science reference|Doyle, S.H., Hubbard, B., Christoffersen, P., Young, T. J., Hofstede, C., Bougamont, M., Box, J. E. & Hubbard, A. 2018. Physical conditions of fast glacier flow: 1. Measurements from boreholes drilled to the bed of Store Glacier, West Greenland, Journal of Geophysical Research: Earth Surface, DOI: 10.1002/2017JF004529.
Science DOI|10.1002/2017JF004529
Date|2014
Longitude [°E]|
Latitude [°N]|
Location source|Doyle, 2018
Depth of top measurement [m]|
Depth of bottom measurement [m]|
Ice thickness [m]|
Coverage [% of thickness]|#DIV/0!
Ice thickness source|
Measured from: Top, Bottom, Relative|
General_Note|
Temperature_note|
Thickness_note|
Location_note|
