Borehole ID|Jakobshavn89A
Place Name|Jakobshavn Isbræ
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|M. Lüthi email
Data DOI|
Science Reference|Iken, A., Echelmeyer, Κ., Harrison, W., Funk, M.: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part I. Measurements of temperature and water level in deep boreholes , Journal of Glaciology 39(131), Cambridge University Press (CUP), 15–25, 1993 
Science DOI|10.3189/S0022143000015689
Date|1989
Longitude [°E]|-48.763000000000005
Latitude [°N]|69.169
Location source|Colgan, 2021
Depth of top measurement [m]|2.0
Depth of bottom measurement [m]|1535.0
Ice thickness [m]|1540
Coverage [% of thickness]|100
Ice thickness source|Iken1993
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
