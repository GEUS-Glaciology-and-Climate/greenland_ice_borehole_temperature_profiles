Borehole ID|td2
Descriptive Name|
Area|Paakitsoq
Data reference|Unknown PDF: See td1
Data DOI|
Science reference|
Science DOI|
Date|1988-05-19
Longitude [°E]|-50.13
Latitude [°N]|69.45
Location source|Unknown PDF: See td1
Depth of top measurement [m]|27.0
Depth of bottom measurement [m]|202.0
Ice thickness [m]|470
Coverage [% of thickness]|37
Ice thickness source|Unknown PDF: See td1
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
