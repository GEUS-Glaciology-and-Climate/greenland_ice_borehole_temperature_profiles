Borehole ID|Jakobshavn89A
Place name|Jakobshavn Isbræ
Geographic location|Central West Greenland
Site type|Ice sheet
Data Source|Lüthi email
Data DOI|
Science Source|Iken, A., Echelmeyer, Κ., Harrison, W., Funk, M.: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part I. Measurements of temperature and water level in deep boreholes , Journal of Glaciology 39(131), Cambridge University Press (CUP), 15–25, 1993 
Science DOI|10.3189/S0022143000015689
Date|1989
Longitude [°E]|-48.763
Latitude [°N]|69.169
Location Source|10.5194/essd-14-2209-2022
Depth of top measurement [m]|2.0
Depth of bottom measurement [m]|1535
Ice thickness [m]|1540
Coverage [% of thickness]|100
Ice thickness source|Iken, 1993
Note|
