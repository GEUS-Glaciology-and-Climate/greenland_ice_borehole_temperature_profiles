Borehole ID|StationCentrale
Place name|Station Centrale
Geographic location|Northwest Greenland
Ice type|Ice sheet
Data Source|Table in science source
Data DOI|
Science Source|Heuberger, J.-C. 1954. Expéditions Polaires Françaises: Missions Paul-Emil Victor. Glaciologie Groenland Volume 1: Forages sur l'inlandsis. Hermann & Cle, Éditeurs. Paris.
Science DOI|
Date|1950
Longitude [°E]|-40.63
Latitude [°N]|70.92
Location Source|https://en.wikipedia.org/wiki/List_of_ice_cores#Greenland
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|150
Ice thickness [m]|3037
Coverage [% of thickness]|5
Ice thickness source|BedMachine_V3
Velocity [m/yr]|14.5
Note|
