Borehole ID|law_2021
Descriptive Name|R30_BH19c
Area|Store Glacier
Data reference|Law, R., Christoffersen, P., Hubbard, B., & Doyle, S. (2021). Distributed temperature sensing data from a borehole drilled to the base of Sermeq Kujalleq (Store Glacier), Greenland, in July 2019 [Dataset]. https://doi.org/10.17863/CAM.65812
Data DOI|10.17863/CAM.65812
Science reference|"Law, Robert, Poul Christoffersen, Bryn Hubbard, Samuel H. Doyle, Thomas R. Chudley, Charlotte M. Schoonman, Marion Bougamont et al. ""Thermodynamics of a fast-moving Greenlandic outlet glacier revealed by fiber-optic distributed temperature sensing."" Science Advances 7, no. 20 (2021): eabe7136."
Science DOI|10.1126/sciadv.abe7136
Date|
Longitude [°E]|-50.09
Latitude [°N]|70.57
Location source|Law (2021)
Depth of top measurement [m]|
Depth of bottom measurement [m]|
Ice thickness [m]|1043
Coverage [% of thickness]|0
Ice thickness source|Law (2021)
Measured from: Top, Bottom, Relative|
General_Note|
Temperature_note|
Thickness_note|
Location_note|
