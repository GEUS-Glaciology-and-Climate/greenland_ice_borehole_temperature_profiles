Borehole ID|Laika_75e
Place name|Laika Ice Cap
Geographic location|Canadian Arctic North
Ice type|Ice cap
Data Source|Graphic in science source
Data DOI|
Science Source|Blatter, Heinz, Kappenberger, Giovanni: Mass Balance and Thermal Regime of Laika Ice Cap, Coburg Island, N.W.T., Canada , Journal of Glaciology 34(116), International Glaciological Society, 102–110, 1988
Science DOI|10.3189/s0022143000009126
Date|1975-08
Longitude [°E]|-79.1801
Latitude [°N]|75.8817
Location Source|10.3189/s0022143000009126
Depth of top measurement [m]|9.0
Depth of bottom measurement [m]|39
Ice thickness [m]|48
Coverage [% of thickness]|63
Ice thickness source|See science reference
Note|Temperature, location, and thickness digitized by M. Jacquemart
