Name|grip
Alternate name|GRIP
Data source|Johnsen, Sigfus J., Dahl-Jensen, Dorthe, Dansgaard, Willi, Gundestrup, Niels: Greenland palaeotemperatures derived from GRIP bore hole temperature and ice core isotope profiles , Tellus B: Chemical and Physical Meteorology 47(5), Informa UK Limited, 624–629, 1 1995 
Drill year(s)|1989-1992 (Vinther, 2008)
Data year(s)|
Longitude [°E]|-37.64
Latitude [°N]|72.58
Approximate location name|
Location source|Vinther (2008)
Ice thickness [m]|3027
Ice thickness year|
Ice thickness source|Montagnat, M., Azuma, N., Dahl-Jensen, D., Eichler, J., Fujita, S., Gillet-Chaulet, F., Kipfstuhl, S., Samyn, D., Svensson, A., Weikusat, I.: Fabric along the NEEM ice core, Greenland, and its comparison with GRIP and NGRIP ice cores , The Cryosphere 8(4), Copernicus GmbH, 1129–1138, 7 2014 
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|107.0
Depth of bottom measurement [m]|3023.0
