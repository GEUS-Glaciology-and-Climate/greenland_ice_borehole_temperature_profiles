Borehole ID|isua_10
Descriptive Name|Isua
Area|
Data reference|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 
Data DOI|
Science reference|
Science DOI|
Date|1972-1973
Longitude [°E]|-49.75
Latitude [°N]|65.2093
Location source|
Depth of top measurement [m]|5.0
Depth of bottom measurement [m]|95.0
Ice thickness [m]|97
Coverage [% of thickness]|93
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
