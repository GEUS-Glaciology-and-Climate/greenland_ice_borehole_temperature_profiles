Borehole ID|dye_3
Descriptive Name|DYE-3
Area|South Greenland
Data reference|Gundestrup, N. S., Hansen, B. Lyle: Bore-Hole Survey at Dye 3, South Greenland , Journal of Glaciology 30(106), Cambridge University Press (CUP), 282–288, 1984 
Data DOI|
Science reference|
Science DOI|
Date|1983
Longitude [°E]|-43.816667
Latitude [°N]|65.18333299999999
Location source|See data source
Depth of top measurement [m]|152.0
Depth of bottom measurement [m]|2030.0
Ice thickness [m]|2038
Coverage [% of thickness]|92
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
