Borehole ID|Isunnguata_27km-11A
Place name|Isunnguata Sermia
Geographic location|Central West Greenland
Site type|Ice sheet
Data Source|Joel Harper and Toby Meierbachtol. 2021. Western Greenland Ice Sheet ice temperature profiles, 2010-2012. Arctic Data Center
Data DOI|10.18739/A2QV3C51Q
Science Source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A945
Date|2011
Longitude [°E]|-49.71952
Latitude [°N]|67.19518
Location Source|T. Meierbachtol email
Depth of top measurement [m]|218.0
Depth of bottom measurement [m]|368
Ice thickness [m]|458
Coverage [% of thickness]|33
Ice thickness source|T. Meierbachtol email
Note|See data in M1-10 folder; Harrington 2015 name: S3-A
