Name|foxx2
Alternate name|FOXX2
Data source|Lüthi, Martin P., Ryser, Claudia, Andrews, Lauren C., Catania, Ginny A., Funk, Martin, Hawley, Robert L., Hoffman, Matthew J., Neumann, Thomas A.: Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming , The Cryosphere 9(1), 245–253, 2015 
Drill year(s)|
Data year(s)|2011-2013
Longitude [°E]|
Latitude [°N]|
Approximate location name|Paakitsoq
Location source|
Ice thickness [m]|
Ice thickness year|
Ice thickness source|
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|8.6
Depth of bottom measurement [m]|285.9
