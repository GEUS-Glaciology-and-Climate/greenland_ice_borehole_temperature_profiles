Borehole ID|Agassiz79a
Place name|Agassiz Ice Cap
Geographic location|Canadian Arctic North
Site type|Ice cap
Data Source|Zdanowicz email
Data DOI|
Science Source|Clarke, G., D. Fisher and E. Waddington. Wind pumping: A potentially significant heat source in ice sheets , The Physical Basis of Ice Sheet Modelling in Proceedings of the Vancouver Symposium, IAHS , volume 170, 169–180, 1987
Science DOI|
Date|1979
Longitude [°E]|-73.1
Latitude [°N]|80.7
Location Source|Vinther, 2008
Depth of top measurement [m]|12.0
Depth of bottom measurement [m]|142
Ice thickness [m]|142
Coverage [% of thickness]|92
Ice thickness source|See data source 
Note|Ice thickness from data does not match ice thickness from Vinther (2008); Location approximate
