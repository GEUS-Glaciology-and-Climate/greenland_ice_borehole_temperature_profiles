Borehole ID|FOXX1
Place name|FOXX
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Graphic in science source
Data DOI|
Science Source|Lüthi, M., C. Ryser, L. Andrews et al. 2015. Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming. The Cryosphere. 9: 245-253. 
Science DOI|10.5194/tc-9-245-2015
Date|2011-2013 @LUTHI
Longitude [°E]|-49.8803
Latitude [°N]|69.4464
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|6.0
Depth of bottom measurement [m]|611
Ice thickness [m]|631
Coverage [% of thickness]|96
Ice thickness source|Martin Luthi
Note|
