Borehole ID|NGRIP
Place Name|NGRIP
Geographic Location|Central Greenland
Ice Type|Ice sheet
Data Reference|G. Clow email
Data DOI|
Science Reference|Buchardt, S. and D. Dahl-Jensen. 2007. Estimating the basal melt rate at NorthGRIP using a Monte Carlo technique. Annals of Glaciology. 45: 137-142. 
Science DOI|10.3189/172756407782282435
Date|2003
Longitude [°E]|-42.32
Latitude [°N]|75.1
Location source|Vinther (2008)
Depth of top measurement [m]|82.0
Depth of bottom measurement [m]|2992
Ice thickness [m]|3085
Coverage [% of thickness]|94
Ice thickness source|See data source email
General_Note|
Temperature_note|
Thickness_note|
Location_note|
