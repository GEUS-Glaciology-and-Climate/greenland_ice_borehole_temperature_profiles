Borehole ID|Penny96
Place Name|Penny Ice Cap
Geographic Location|Canadian Arctic South
Ice Type|Ice cap
Data Reference|W. Colgan email
Data DOI|
Science Reference|Fisher, D., R. Koerner, J. Bourgeois et al. 1998. Penny Ice Cap Cores, Baffin Island, Canada, and the Wisconsinan Foxe Dome Connection: Two States of Hudson Bay Ice Cover. Science. 279: 692-695. 
Science DOI|10.1126/science.279.5351.692
Date|1996
Longitude [°E]|-65.2
Latitude [°N]|67.3
Location source|Colgan, 2021
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|176.0
Ice thickness [m]|176
Coverage [% of thickness]|94
Ice thickness source|Data file + WIC email (see also Fisher 1998)
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
