Borehole ID|Tuto_D-11
Place name|Tuto Ramp
Geographic location|Northwest Greenland
Site type|Ice sheet
Data Source|Graphic in science source
Data DOI|
Science Source|Davis, RM: Approach roads, Greenland 1960–1964 , Technical Report 133. Corps of Engineers, Cold Regions Research & Engineering Laboratory , 1967 
Science DOI|
Date|1962-08-15
Longitude [°E]|-68.2873
Latitude [°N]|76.4113
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|0.0
Depth of bottom measurement [m]|48
Ice thickness [m]|48
Coverage [% of thickness]|100
Ice thickness source|See data source
Note|
