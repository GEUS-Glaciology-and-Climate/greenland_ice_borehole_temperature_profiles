Borehole ID|TD1_88
Place Name|Paakitsoq
Geographic Location|Central West Greenland
Ice Type|
Data Reference|Unknown PDF: Shallow88II.pdf
Data DOI|
Science Reference|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1988-05-19
Longitude [°E]|-50.13
Latitude [°N]|69.45
Location source|Colgan2021
Depth of top measurement [m]|50.0
Depth of bottom measurement [m]|300.0
Ice thickness [m]|300.0
Coverage [% of thickness]|83
Ice thickness source|Unknown PDF: Shallow88II.pdf
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
