Borehole ID|FladeIsblink06
Place name|Flade Isblink Ice Cap
Geographic location|Northeast Greenland
Site type|Ice cap
Data Source|Dalh-Jensen email
Data DOI|
Science Source|Lemark, A. and D. Dahl-Jensen. 2010. A study of the Flade Isblink ice cap using a simple ice flow model. Master's thesis. Niels Bohr Institute, Copenhagen University.
Science DOI|
Date|2006
Longitude [°E]|-15.7029
Latitude [°N]|81.2926
Location Source|10.5194/essd-14-2209-2022
Depth of top measurement [m]|80.0
Depth of bottom measurement [m]|420
Ice thickness [m]|540
Coverage [% of thickness]|63
Ice thickness source|W. Colgan email
Note|
