Name|isua_11
Alternate name|Isua
Data source|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 
Drill year(s)|
Data year(s)|1972-1973
Longitude [°E]|-49.7510
Latitude [°N]|65.2072
Approximate location name|
Location source|
Ice thickness [m]|120
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|25.0
Depth of bottom measurement [m]|116.0
