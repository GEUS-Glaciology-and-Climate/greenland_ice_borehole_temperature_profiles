Borehole ID|PrinceWales05
Place name|Prince of Wales Ice Cap
Geographic location|Canadian Arctic North
Site type|Ice cap
Data Source|Zdanowicz email
Data DOI|
Science Source|Kinnard, C., R. Koerner, C. Zdanowicz et al. 2008. Stratigraphic analysis of an ice core from the Prince of Wales Icefield, Ellesmere Island, Arctic Canada, using digital image analysis: High‐resolution density, past summer warmth reconstruction, and melt effect on ice core solid conductivity. Journal of Geophysical Research. 113: D24120. 
Science DOI|10.1029/2008JD011083
Date|2005-05-15
Longitude [°E]|-80.395
Latitude [°N]|78.3897
Location Source|10.5194/essd-14-2209-2022
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|176
Ice thickness [m]|176
Coverage [% of thickness]|94
Ice thickness source|W. Colgan email
Note|
