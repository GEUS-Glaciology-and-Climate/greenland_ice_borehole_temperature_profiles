Borehole ID|GISP2
Place Name|GISP2
Geographic Location|Central Greenland
Ice Type|Ice sheet
Data Reference|G. Clow email
Data DOI|
Science Reference|MacGregor, J., J. Li, J. Paden et al. 2015. Radar attenuation and temperature within the Greenland Ice Sheet. Journal of Geophysical Research. 120: 983-1008. 
Science DOI|10.1002/2014JF003418
Date|1996-06-02
Longitude [°E]|-38.4667
Latitude [°N]|72.5833
Location source|Colgan, 2021
Depth of top measurement [m]|73.0
Depth of bottom measurement [m]|3053.0
Ice thickness [m]|3100
Coverage [% of thickness]|96
Ice thickness source|Hodge 1990?
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|Location from Geothermal Database
