Borehole ID|CampCentury
Place name|Camp Century
Geographic location|Northwest Greenland
Ice type|Ice cap
Data Source|Graphic in science source
Data DOI|
Science Source|Weertman, J.: Comparison between measured and theoretical temperature profiles of the Camp Century, Greenland, Borehole , Journal of Geophysical Research 73(8), American Geophysical Union (AGU), 2691–2700, 4 1968
Science DOI|10.1029/jb073i008p02691
Date|1966
Longitude [°E]|-61.1097
Latitude [°N]|77.1797
Location Source|Colgan, 2021
Depth of top measurement [m]|9.0
Depth of bottom measurement [m]|1387
Ice thickness [m]|1387
Coverage [% of thickness]|99
Ice thickness source|Weertman1968
Note|
