Borehole ID|Isunnguata_M2-10B
Place name|Isunnguata Sermia
Geographic location|Central West Greenland
Site type|Ice sheet
Data Source|Joel Harper and Toby Meierbachtol. 2021. Western Greenland Ice Sheet ice temperature profiles, 2010-2012. Arctic Data Center
Data DOI|10.18739/A2QV3C51Q
Science Source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A940
Date|2010
Longitude [°E]|-50.06633
Latitude [°N]|67.16704
Location Source|T. Meierbachtol email
Depth of top measurement [m]|6.0
Depth of bottom measurement [m]|131
Ice thickness [m]|146
Coverage [% of thickness]|86
Ice thickness source|T. Meierbachtol email
Note|See data in M1-10 folder; Harrington 2015 name: S1-B
