Borehole ID|Isunnguata_27km-11A
Place name|Isunnguata Sermia
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Meierbachtol email
Data DOI|
Science Source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A942
Date|2011
Longitude [°E]|-49.71952
Latitude [°N]|67.19518000000001
Location Source|Meierbachtol email
Depth of top measurement [m]|218.0
Depth of bottom measurement [m]|368
Ice thickness [m]|458
Coverage [% of thickness]|33
Ice thickness source|T. Meierbachtol email
Note|See data in M1-10 folder; Harrington 2015 name: S3-A
