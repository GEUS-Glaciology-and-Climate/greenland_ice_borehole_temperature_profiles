Borehole ID|GULL5
Place name|Sermeq Avannerleq
Geographic location|Central West Greenland
Site type|Ice sheet
Data Source|Lüthi email
Data DOI|
Science Source|Ryser, C., Lüthi, M. P., Andrews, L. C., Hoffman, M. J., Catania, G. A., Hawley, R. L., ... & Kristensen, S. S. (2014). Sustained high basal motion of the Greenland ice sheet revealed by borehole deformation. Journal of Glaciology, 60(222), 647-660.
Science DOI|10.3189/2014JoG13J196
Date|2011-07-29
Longitude [°E]|-49.7182
Latitude [°N]|69.4524
Location Source|10.3189/2014JoG13J196
Depth of top measurement [m]|307.0
Depth of bottom measurement [m]|707
Ice thickness [m]|707
Coverage [% of thickness]|57
Ice thickness source|Ryser, 2014 (Table 3). 705/707 for thickness
Note|See FOXX1/temperature_foxx_gull_streamlined.org
