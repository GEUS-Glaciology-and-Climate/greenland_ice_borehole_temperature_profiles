Borehole ID|HansTausen_Dome
Place Name|Hans Tausen Dome
Geographic Location|North Greenland
Ice Type|
Data Reference|H. Zekollari email
Data DOI|
Science Reference|Zekollari, Harry, Huybrechts, Philippe, Noël, Brice, van de Berg, Willem Jan, van den Broeke, Michiel R.: Sensitivity, stability and future evolution of the world’s northernmost ice cap, Hans Tausen Iskappe (Greenland) , The Cryosphere 11(2), Copernicus GmbH, 805–825, 3 2017 
Science DOI|10.5194/tc-11-805-2017
Date|1995
Longitude [°E]|-37.47
Latitude [°N]|82.51
Location source|Colgan2021
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|345.0
Ice thickness [m]|345.0
Coverage [% of thickness]|97
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|Only two data points - 10 m and 345 m. Drill date: 10.34194/bullggu.v172.6749 
Temperature_note|
Thickness_note|
Location_note|
