Borehole ID|CampIII_78
Place name|Nunap Kigdlinga
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Table in science source
Data DOI|
Science Source|Stauffer, B., and H. Oeschger. 1979. Temperaturprofile in bohrloechern am rande des Groenlaendischen Inlandeises. Hydrologie und Glaziologie an der ETH Zurich. Mitteilung Nr. 41.
Science DOI|
Date|1978
Longitude [°E]|-49.8
Latitude [°N]|69.722
Location Source|EGIG_CarteNo7
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|90
Ice thickness [m]|539
Coverage [% of thickness]|15
Ice thickness source|BedMachine_V3
Note|See also shallow profiles at boreholes I and III
