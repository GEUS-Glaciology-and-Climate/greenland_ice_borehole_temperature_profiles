Borehole ID|gisp2
Descriptive Name|GISP2, GISP II
Area|
Data reference|G. Clow email
Data DOI|
Science reference|
Science DOI|
Date|1996-06-02
Longitude [°E]|-38.4667
Latitude [°N]|72.5833
Location source|
Depth of top measurement [m]|72.61
Depth of bottom measurement [m]|3053.15
Ice thickness [m]|3100
Coverage [% of thickness]|96
Ice thickness source|Hodge 1990?
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|Location from Geothermal Database
