Borehole ID|tuto_ramp
Descriptive Name|Tuto Ramp
Area|Thule Approach Road(?)
Data reference|Davis, RM: Approach roads, Greenland 1960–1964 , Technical Report 133. Corps of Engineers, Cold Regions Research & Engineering Laboratory , 1967 
Data DOI|
Science reference|
Science DOI|
Date|1962 (August)
Longitude [°E]|-68.287295
Latitude [°N]|76.41133
Location source|
Depth of top measurement [m]|
Depth of bottom measurement [m]|
Ice thickness [m]|48
Coverage [% of thickness]|0
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T(ish)
General_Note|
Temperature_note|
Thickness_note|
Location_note|
