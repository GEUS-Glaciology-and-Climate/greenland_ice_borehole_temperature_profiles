Borehole ID|devon_00
Descriptive Name|Devon borehole
Area|Devon Ice Cap
Data reference|W. Colgan email
Data DOI|
Science reference|
Science DOI|
Date|2000-04-15
Longitude [°E]|-82.14
Latitude [°N]|75.34
Location source|
Depth of top measurement [m]|13.0
Depth of bottom measurement [m]|218.0
Ice thickness [m]|300.55
Coverage [% of thickness]|68
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
