Borehole ID|StationCentrale
Place Name|Station Centrale
Geographic Location|
Ice Type|
Data Reference|
Data DOI|
Science Reference|Heuberger, J.-C. 1954. Expéditions Polaires Françaises: Missions Paul-Emil Victor. Glaciologie Groenland Volume 1: Forages sur l'inlandsis. Hermann & Cle, Éditeurs. Paris.
Science DOI|
Date|
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|150.0
Ice thickness [m]|
Coverage [% of thickness]|
Ice thickness source|
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/files/7082104/heuberger_1954.pdf
Thickness_note|
Location_note|
