Borehole ID|jakobshavn_center
Descriptive Name|
Area|
Data reference|Iken, A., Echelmeyer, Κ., Harrison, W., Funk, M.: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part I. Measurements of temperature and water level in deep boreholes , Journal of Glaciology 39(131), Cambridge University Press (CUP), 15–25, 1993 
Data DOI|
Science reference|
Science DOI|
Date|
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|12.0
Depth of bottom measurement [m]|2410.0
Ice thickness [m]|2495
Coverage [% of thickness]|96
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
