Borehole ID|NGRIP
Place name|NGRIP
Geographic location|Central Greenland
Ice type|Ice sheet
Data Source|Clow email
Data DOI|
Science Source|Buchardt, S. and D. Dahl-Jensen. 2007. Estimating the basal melt rate at NorthGRIP using a Monte Carlo technique. Annals of Glaciology. 45: 137-142. 
Science DOI|10.3189/172756407782282435
Date|2003
Longitude [°E]|-42.32
Latitude [°N]|75.1
Location Source|Vinther, 2008
Depth of top measurement [m]|82.0
Depth of bottom measurement [m]|2992
Ice thickness [m]|3085
Coverage [% of thickness]|94
Ice thickness source|See data source email
Note|
