Borehole ID|Tuto_D-11
Place Name|Tuto Ramp
Geographic Location|Northwest Greenland
Ice Type|
Data Reference|Davis, RM: Approach roads, Greenland 1960–1964 , Technical Report 133. Corps of Engineers, Cold Regions Research & Engineering Laboratory , 1967 
Data DOI|
Science Reference|Davis, RM: Approach roads, Greenland 1960–1964 , Technical Report 133. Corps of Engineers, Cold Regions Research & Engineering Laboratory , 1967 
Science DOI|
Date|1962-08-15
Longitude [°E]|-68.2873
Latitude [°N]|76.4113
Location source|Colgan2021
Depth of top measurement [m]|0.0
Depth of bottom measurement [m]|48.0
Ice thickness [m]|48.0
Coverage [% of thickness]|100
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T(ish)
General_Note|
Temperature_note|
Thickness_note|
Location_note|
