Borehole ID|TD4_91b
Place name|Paakitsoq
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Lüthi email
Data DOI|
Science Source|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1991-08-28
Longitude [°E]|-49.68
Latitude [°N]|69.53
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|3.0
Depth of bottom measurement [m]|493
Ice thickness [m]|660
Coverage [% of thickness]|74
Ice thickness source|Estimate from Martin Luthi
Note|
