Borehole ID|Isunnguata_27km-12A
Place Name|Isunnguata Sermia
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|T. Meierbachtol email
Data DOI|
Science Reference|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A945
Date|2012
Longitude [°E]|-49.71793
Latitude [°N]|67.20421999999999
Location source|T. Meierbachtol email
Depth of top measurement [m]|11.0
Depth of bottom measurement [m]|690.0
Ice thickness [m]|696
Coverage [% of thickness]|98
Ice thickness source|T. Meierbachtol email
Measured from: Top, Bottom, Relative|T
General_Note|See data in M1-10 folder
Temperature_note|
Thickness_note|
Location_note|Harrington 2015 name: S4-A
