Name|meighen
Alternate name|Meighen Ice Cap
Data source|Paterson, W. S. B.: A temperature profile through the Meighen ice cap, Arctic Canada , International Association of Scientific Hydrology 79, 440–449, 1968 
Drill year(s)|
Data year(s)|1965
Longitude [°E]|
Latitude [°N]|
Approximate location name|
Location source|
Ice thickness [m]|121.2
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|1.0
Depth of bottom measurement [m]|121.0
