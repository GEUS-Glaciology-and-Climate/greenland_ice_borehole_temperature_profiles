Borehole ID|hanstausen_hare
Descriptive Name|Hans Tausen Hare
Area|Hans Tausen Ice Cap
Data reference|H. Zekollari email
Data DOI|
Science reference|Zekollari, Harry, Huybrechts, Philippe, Noël, Brice, van de Berg, Willem Jan, van den Broeke, Michiel R.: Sensitivity, stability and future evolution of the world’s northernmost ice cap, Hans Tausen Iskappe (Greenland) , The Cryosphere 11(2), Copernicus GmbH, 805–825, 3 2017 
Science DOI|10.5194/tc-11-805-2017
Date|1995
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|9.0
Depth of bottom measurement [m]|288.0
Ice thickness [m]|289
Coverage [% of thickness]|97
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|Drill date: 10.34194/bullggu.v172.6749 
Temperature_note|
Thickness_note|
Location_note|
