Name|td1
Alternate name|
Data source|Unknown PDF: Shallow88II.pdf
Drill year(s)|
Data year(s)|1988-05-19
Longitude [°E]|-50.13
Latitude [°N]|69.45
Approximate location name|Paakitsoq
Location source|Unknown PDF: Shallow88II.pdf
Ice thickness [m]|300
Ice thickness year|
Ice thickness source|Unknown PDF: Shallow88II.pdf
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|50.0
Depth of bottom measurement [m]|300.0
