Borehole ID|TD5_90
Place name|Paakitsoq
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Lüthi email
Data DOI|
Science Source|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1990-06-09
Longitude [°E]|-49.3
Latitude [°N]|69.57
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|5.0
Depth of bottom measurement [m]|600
Ice thickness [m]|1223
Coverage [% of thickness]|49
Ice thickness source|BedMachine_V3
Note|
