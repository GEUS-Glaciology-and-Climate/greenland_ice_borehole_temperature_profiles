Borehole ID|jakobshavn_sheet
Descriptive Name|
Area|
Data reference|Lüthi, Martin, Funk, Martin, Iken, Almut, Gogineni, Shivaprasad, Truffer, Martin: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part III. Measurements of ice deformation, temperature and cross-borehole conductivity in boreholes to the bedrock , Journal of Glaciology 48(162), 369–385, 2002 
Data DOI|
Science reference|
Science DOI|
Date|1995
Longitude [°E]|-48.68713
Latitude [°N]|69.235046
Location source|See data source
Depth of top measurement [m]|19.0
Depth of bottom measurement [m]|798.0
Ice thickness [m]|828
Coverage [% of thickness]|94
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|Location from Geothermal Database
