Name|ngrip
Alternate name|NGRIP
Data source|G. Clow email
Drill year(s)|1996-2004 (Vinther, 2008)
Data year(s)|
Longitude [°E]|-42.32
Latitude [°N]|75.10
Approximate location name|
Location source|Vinther (2008)
Ice thickness [m]|3085
Ice thickness year|
Ice thickness source|See data source email
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|81.89
Depth of bottom measurement [m]|2992.47
