Name|template
Alternate name|Template Borehole
Data source|Reference
Data year(s)|YYYY
Depth of top measurement [m]|float
Depth of bottom measurement [m]|float
Drill year(s)|YYYY
Longitude [°E]|decimal degree
Latitude [°N]|decimal degree
Approximate location name|Location Name
Location source|Reference
Ice thickness [m]|float
Ice thickness year|YYYY
Ice thickness source|Reference
Surface velocity [m yr^-1]|float
Surface velocity year|YYYY
Surface velocity source|Reference
Measured from: Top, Bottom, Relative|T/B/R
