Borehole ID|Store_R30_BH19c
Place Name|Store Glacier
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|R. Law email
Data DOI|
Science Reference|"Law, Robert, Poul Christoffersen, Bryn Hubbard, Samuel H. Doyle, Thomas R. Chudley, Charlotte M. Schoonman, Marion Bougamont et al. ""Thermodynamics of a fast-moving Greenlandic outlet glacier revealed by fiber-optic distributed temperature sensing."" Science Advances 7, no. 20 (2021): eabe7136."
Science DOI|10.1126/sciadv.abe7136
Date|2019-08-13
Longitude [°E]|-50.09
Latitude [°N]|70.57
Location source|Law (2021)
Depth of top measurement [m]|0.09
Depth of bottom measurement [m]|1044
Ice thickness [m]|1044
Coverage [% of thickness]|100
Ice thickness source|Law (2021)
General_Note|See also: 10.5285/ecf81955-b829-4f91-ae90-b9bc947f8c60
Temperature_note|
Thickness_note|
Location_note|
