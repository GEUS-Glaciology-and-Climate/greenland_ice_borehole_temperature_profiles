Name|gisp2
Alternate name|GISP2; GISP II
Data source|Cuffey, Kurt M., Alley, Richard B., Grootes, Pieter M., Anandakrishnan, Sridhar: Toward using borehole temperatures to calibrate an isotopic paleothermometer in central Greenland , Palaeogeography, Palaeoclimatology, Palaeoecology 98(2-4), Elsevier BV, 265–268, 12 1992 
Drill year(s)|
Data year(s)|1989,1990
Longitude [°E]|
Latitude [°N]|
Approximate location name|Russell / Leverett ?
Location source|
Ice thickness [m]|3100
Ice thickness year|
Ice thickness source|Hodge 1990?
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|37.0
Depth of bottom measurement [m]|216.0
