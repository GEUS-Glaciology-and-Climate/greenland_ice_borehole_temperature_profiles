Borehole ID|harrington_2015_27km-12C
Descriptive Name|27km-12C
Area|
Data reference|T. Meierbachtol email
Data DOI|
Science reference|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A947
Date|2012
Longitude [°E]|-49.718114
Latitude [°N]|67.20382
Location source|T. Meierbachtol email
Depth of top measurement [m]|17.0
Depth of bottom measurement [m]|688.0
Ice thickness [m]|696
Coverage [% of thickness]|96
Ice thickness source|T. Meierbachtol email
Measured from: Top, Bottom, Relative|T
General_Note|See data in M1-10 folder
Temperature_note|
Thickness_note|
Location_note|Harrington 2015 name: S4-C
