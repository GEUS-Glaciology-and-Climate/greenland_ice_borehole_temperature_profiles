Borehole ID|TD5_91
Place Name|Paakitsoq
Geographic Location|Central West Greenland
Ice Type|
Data Reference|Unknown PDF: See td1 and Lüthi (2015)
Data DOI|
Science Reference|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1991-05-25
Longitude [°E]|-49.3
Latitude [°N]|69.57
Location source|Colgan2021
Depth of top measurement [m]|5.0
Depth of bottom measurement [m]|600.0
Ice thickness [m]|1223.0
Coverage [% of thickness]|49
Ice thickness source|BedMachine_V3
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
