Borehole ID|CampIII_78b
Place Name|Nunap Kigdlinga
Geographic Location|
Ice Type|
Data Reference|Stauffer, 1979
Data DOI|
Science Reference|
Science DOI|
Date|1978
Longitude [°E]|-50.0917
Latitude [°N]|69.7176
Location source|M. Lüthi email
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|90
Ice thickness [m]|
Coverage [% of thickness]|#DIV/0!
Ice thickness source|
General_Note|See also shallow profiles at boreholes I and III
Temperature_note|Digitized from https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/files/7185440/stauffer_1979.pdf
Thickness_note|
Location_note|
