Name|ngrip
Alternate name|NGRIP
Data source|Dahl-Jensen, Dorthe, Gundestrup, Niels, Gogineni, S Prasad, Miller, Heinz: Basal melt at NorthGRIP modeled from borehole, ice-core and radio-echo sounder observations , Annals of Glaciology 37, International Glaciological Society, 207–212, 2003 
Drill year(s)|1996-2004 (Vinther, 2008)
Data year(s)|
Longitude [°E]|-42.32
Latitude [°N]|75.10
Approximate location name|
Location source|Vinther (2008)
Ice thickness [m]|3080
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|204.0
Depth of bottom measurement [m]|2888.0
