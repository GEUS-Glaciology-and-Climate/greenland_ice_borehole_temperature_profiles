Borehole ID|camp_vi
Descriptive Name|Camp VI
Area|
Data reference|Digitization from published graphic
Data DOI|
Science reference|
Science DOI|
Date|1950?
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|4.0
Depth of bottom measurement [m]|125.0
Ice thickness [m]|
Coverage [% of thickness]|#DIV/0!
Ice thickness source|
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
