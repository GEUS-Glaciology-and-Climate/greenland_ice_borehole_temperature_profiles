Borehole ID|gull
Descriptive Name|GULL
Area|Paakitsoq
Data reference|Lüthi, Martin P., Ryser, Claudia, Andrews, Lauren C., Catania, Ginny A., Funk, Martin, Hawley, Robert L., Hoffman, Matthew J., Neumann, Thomas A.: Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming , The Cryosphere 9(1), 245–253, 2015 
Data DOI|
Science reference|
Science DOI|
Date|2011-2013
Longitude [°E]|-49.7142167
Latitude [°N]|69.4526
Location source|
Depth of top measurement [m]|4.0
Depth of bottom measurement [m]|704.0
Ice thickness [m]|703
Coverage [% of thickness]|100
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|Location from Geothermal Database
