Borehole ID|Store_S30
Place Name|Store Glacier
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|Doyle, Samuel; Hubbard, Bryn; Christoffersen, Poul; Young, Tun Jan; Hofstede, Coen; Bougamont, Marion; et al. (2018): SAFIRE borehole, AWS and GPS datasets. figshare. Dataset. https://doi.org/10.6084/m9.figshare.5745294.v1 
Data DOI|10.6084/m9.figshare.5745294.v1
Science Reference|Doyle, S.H., Hubbard, B., Christoffersen, P., Young, T. J., Hofstede, C., Bougamont, M., Box, J. E. & Hubbard, A. 2018. Physical conditions of fast glacier flow: 1. Measurements from boreholes drilled to the bed of Store Glacier, West Greenland, Journal of Geophysical Research: Earth Surface, DOI: 10.1002/2017JF004529.
Science DOI|10.1002/2017JF004529
Date|2014
Longitude [°E]|-49.9167
Latitude [°N]|70.5167
Location source|Doyle, 2018
Depth of top measurement [m]|102.0
Depth of bottom measurement [m]|604
Ice thickness [m]|600
Coverage [% of thickness]|84
Ice thickness source|Doyle (2018)
General_Note|
Temperature_note|
Thickness_note|
Location_note|
