Borehole ID|GRIP
Place name|GRIP
Geographic location|Central Greenland
Ice type|Ice sheet
Data Source|Clow email
Data DOI|
Science Source|MacGregor, J., J. Li, J. Paden et al. 2015. Radar attenuation and temperature within the Greenland Ice Sheet. Journal of Geophysical Research. 120: 983-1008. 
Science DOI|10.1002/2014JF003418
Date|1998
Longitude [°E]|-37.64
Latitude [°N]|72.58
Location Source|Vinther, 2008
Depth of top measurement [m]|41.0
Depth of bottom measurement [m]|3029
Ice thickness [m]|3029
Coverage [% of thickness]|99
Ice thickness source|G. Clow email
Note|
