Name|flade_isblink
Alternate name|Flade Isblink
Data source|Dorthe Dalh-Jensen (personal comm.)
Drill year(s)|
Data year(s)|
Longitude [°E]|-15.7029
Latitude [°N]|81.2926
Approximate location name|
Location source|
Ice thickness [m]|540
Ice thickness year|
Ice thickness source|See WIC email
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|80.0
Depth of bottom measurement [m]|420.0
