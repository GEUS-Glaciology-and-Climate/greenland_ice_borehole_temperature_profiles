Borehole ID|FladeIsblink06
Place Name|Flade Isblink Ice Cap
Geographic Location|Northeast Greenland
Ice Type|Ice cap
Data Reference|D. Dalh-Jensen email
Data DOI|
Science Reference|Lemark, A. and D. Dahl-Jensen. 2010. A study of the Flade Isblink ice cap using a simple ice flow model. Master's thesis. Niels Bohr Institute, Copenhagen University.
Science DOI|
Date|2006
Longitude [°E]|-15.7029
Latitude [°N]|81.2926
Location source|Colgan, 2021
Depth of top measurement [m]|80.0
Depth of bottom measurement [m]|420
Ice thickness [m]|540
Coverage [% of thickness]|63
Ice thickness source|See WIC email
General_Note|
Temperature_note|
Thickness_note|
Location_note|
