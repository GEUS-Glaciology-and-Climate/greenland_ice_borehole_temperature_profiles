Borehole ID|HansTausen_Dome
Place name|Hans Tausen Dome
Geographic location|North Greenland
Site type|Ice cap
Data Source|E. Zwelty, Issue #50, and Reeh, Niels, ed. Report on Activities and Results 1993-1995 for Hans Tavsen Ice Cap Project: Glacier and Climate Change Research, North Greenland. 1995. Fig. 6.
Data DOI|
Science Source|Zekollari, Harry, Huybrechts, Philippe, Noël, Brice, van de Berg, Willem Jan, van den Broeke, Michiel R.: Sensitivity, stability and future evolution of the world’s northernmost ice cap, Hans Tausen Iskappe (Greenland) , The Cryosphere 11(2), Copernicus GmbH, 805–825, 3 2017 
Science DOI|10.5194/tc-11-805-2017
Date|1995
Longitude [°E]|-37.47
Latitude [°N]|82.51
Location Source|10.5194/essd-14-2209-2022
Depth of top measurement [m]|12.0
Depth of bottom measurement [m]|341
Ice thickness [m]|345
Coverage [% of thickness]|95
Ice thickness source|See data source
Note|Drill date: 10.34194/bullggu.v172.6749 
