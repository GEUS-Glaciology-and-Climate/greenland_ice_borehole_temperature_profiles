Borehole ID|Store_R30_BH19c
Place name|Store Glacier
Geographic location|Central West Greenland
Site type|Ice sheet
Data Source|Law email
Data DOI|
Science Source|"Law, Robert, Poul Christoffersen, Bryn Hubbard, Samuel H. Doyle, Thomas R. Chudley, Charlotte M. Schoonman, Marion Bougamont et al. ""Thermodynamics of a fast-moving Greenlandic outlet glacier revealed by fiber-optic distributed temperature sensing."" Science Advances 7, no. 20 (2021): eabe7136."
Science DOI|10.1126/sciadv.abe7136
Date|2019-08-13
Longitude [°E]|-50.09
Latitude [°N]|70.57
Location Source|Law, 2021
Depth of top measurement [m]|0.09
Depth of bottom measurement [m]|1044
Ice thickness [m]|1044
Coverage [% of thickness]|100
Ice thickness source|Law (2021)
Note|See also: 10.5285/ecf81955-b829-4f91-ae90-b9bc947f8c60 (Note, both fibre optic DTS and thermistor data are presented in Law et al. (2021))
