Borehole ID|h2015_s2a
Descriptive Name|13km_S2A
Area|
Data reference|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Data DOI|
Science reference|
Science DOI|
Date|2010
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|3.5
Depth of bottom measurement [m]|559.0
Ice thickness [m]|
Coverage [% of thickness]|#DIV/0!
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
