Name|devon_72
Alternate name|Devon borehole
Data source|Paterson, W. S. B., Clarke, G. K. C.: Comparison of theoretical and observed temperature profiles in Devon Island ice cap, Canada , Geophysical Journal International 55(3), Oxford University Press (OUP), 615–632, 12 1978 
Drill year(s)|
Data year(s)|
Longitude [°E]|-82.14
Latitude [°N]|75.34
Approximate location name|Devon Ice Cap
Location source|
Ice thickness [m]|299
Ice thickness year|drill year
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|9
Depth of bottom measurement [m]|299
