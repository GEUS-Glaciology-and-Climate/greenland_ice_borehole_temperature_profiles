Borehole ID|Barnes_T0975_1976
Place name|Barnes Ice Cap
Geographic location|Canadian Arctic South
Ice type|Ice cap
Data Source|Graphic in science source
Data DOI|
Science Source|Hooke, Roger LeB., Alexander, E. Calvin, Gustafson, Robert J.: Temperature profiles in the Barnes Ice Cap, Baffin Island, Canada, and heat flux from the subglacial terrane , Canadian Journal of Earth Sciences 17(9), Canadian Science Publishing, 1174–1188, sep 1980
Science DOI|10.1139/e80-124
Date|1976-06-22
Longitude [°E]|-72.1103
Latitude [°N]|69.79795
Location Source|Location digitized by M. Jacquemart from Gilbert (2016)
Depth of top measurement [m]|0.0
Depth of bottom measurement [m]|47
Ice thickness [m]|115
Coverage [% of thickness]|41
Ice thickness source|See science source
Note|"Date is ""Date completed"" from Hooke (1980) Table 1 Column 2 + Days to final measurement (Column 3); Temperature and location digitized by M. Jacquemart from Gilbert (2016)"
