Name|camp_century
Alternate name|Camp Century
Data source|Weertman, J.: Comparison betwe
Drill year(s)|nan
Data year(s)|nan
Longitude [°E]|nan
Latitude [°N]|nan
Approximate location name|Camp Century
Location source|?
Ice thickness [m]|1387
Ice thickness year|?
Ice thickness source|?
Surface velocity [m yr^-1]|nan
Surface velocity year|nan
Surface velocity source|nan
Measured from: Top, Bottom, Relative|B
Depth of top measurement [m]|9.0
Depth of bottom measurement [m]|1387.0
Coverage [% of thickness]|99
