Borehole ID|Barnes_24.55_T_1975
Place name|Barnes Ice Cap
Geographic location|Canadian Arctic South
Site type|Ice cap
Data Source|Table in science source
Data DOI|
Science Source|Classen, D. F.: Temperature profiles for the Barnes Ice Cap surge zone , Journal of Glaciology 18(80), International Glaciological Society, 391–405, 1977
Science DOI|10.3189/s0022143000021079
Date|1975-07-02
Longitude [°E]|-72.1104
Latitude [°N]|69.54665509
Location Source|Location digitized by M. Jacquemart from Classen (1977) and modern aerial images
Depth of top measurement [m]|28.0
Depth of bottom measurement [m]|88
Ice thickness [m]|115
Coverage [% of thickness]|52
Ice thickness source|See science source
Note|Location digitized by M. Jacquemart
