Name|site_ii
Alternate name|Site II
Data source|Hansen, B. L., Landauer, J. K.: Some results of ice cap drill hole measurements, Union Geodesique et Geophysique Internationale. Association Internationale d'Hydrologie Scientifique 47, 313–317, 1958 
Drill year(s)|1957 (Summer)
Data year(s)|1958 (late June)
Longitude [°E]|-56.066667
Latitude [°N]|76.983333
Approximate location name|
Location source|WIC Email
Ice thickness [m]|1851
Ice thickness year|
Ice thickness source|BedMachine
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|
Depth of bottom measurement [m]|
