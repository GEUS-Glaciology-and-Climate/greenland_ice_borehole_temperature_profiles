Borehole ID|Renland88
Place Name|Renland Ice Cap
Geographic Location|Central East Greenland
Ice Type|Ice cap
Data Reference|B. M. Vinther email
Data DOI|
Science Reference|Hansson, M. 1994. The Renland ice core. A Northern Hemisphere record of aerosol composition over 120,000 years. Tellus B. 46: 390-418.
Science DOI|10.3402/tellusb.v46i5.15813
Date|1988
Longitude [°E]|-26.768
Latitude [°N]|71.306
Location source|Email and Vinther (2008)
Depth of top measurement [m]|15.0
Depth of bottom measurement [m]|300.0
Ice thickness [m]|324
Coverage [% of thickness]|88
Ice thickness source|Vinther, B. M., Clausen, H. B., Fisher, D. A., Koerner, R. M., Johnsen, S. J., Andersen, K. K., Dahl-Jensen, D., Rasmussen, S. O., Steffensen, J. P., Svensson, A. M.: Synchronizing ice cores from the Renland and Agassiz ice caps to the Greenland Ice Core Chronology , Journal of Geophysical Research 113(D8), American Geophysical Union (AGU), 4 2008 
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
