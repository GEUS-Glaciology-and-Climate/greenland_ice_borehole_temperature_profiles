Borehole ID|Isua_11
Place Name|Isua
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 
Data DOI|
Science Reference|Colebeck, S. and A. Gow. 1979. The margin of the Greenland Ice Sheet at Isua. Journal of Glaciology. 24: 155-165. 
Science DOI|10.3189/S0022143000014714
Date|1972-1973
Longitude [°E]|-49.751000000000005
Latitude [°N]|65.2072
Location source|Colgan, 2021
Depth of top measurement [m]|25.0
Depth of bottom measurement [m]|116
Ice thickness [m]|120
Coverage [% of thickness]|76
Ice thickness source|See data source
General_Note|
Temperature_note|Digitized from graphic
Thickness_note|
Location_note|
