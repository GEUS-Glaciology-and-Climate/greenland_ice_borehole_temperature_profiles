Borehole ID|isua_14
Descriptive Name|Isua
Area|
Data reference|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 
Data DOI|
Science reference|
Science DOI|
Date|1972-1973
Longitude [°E]|-49.7443
Latitude [°N]|65.2058
Location source|
Depth of top measurement [m]|6.0
Depth of bottom measurement [m]|237.0
Ice thickness [m]|299
Coverage [% of thickness]|77
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
