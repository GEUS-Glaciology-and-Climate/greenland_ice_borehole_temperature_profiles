Borehole ID|SiteII
Place Name|Site II
Geographic Location|Northwest Greenland
Ice Type|
Data Reference|Hansen, B. L., Landauer, J. K.: Some results of ice cap drill hole measurements, Union Geodesique et Geophysique Internationale. Association Internationale d'Hydrologie Scientifique 47, 313–317, 1958 
Data DOI|
Science Reference|Hansen, B. and J. Landauer. 1958. Some results of ice cap drill hole measurements. IASH Publication. 47: 313-317.
Science DOI|
Date|1958-06-25
Longitude [°E]|-56.07
Latitude [°N]|76.98
Location source|Colgan2021
Depth of top measurement [m]|16.0
Depth of bottom measurement [m]|410.0
Ice thickness [m]|1851.0
Coverage [% of thickness]|21
Ice thickness source|BedMachine_V3
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
