Borehole ID|CVI_EPF
Place Name|Camp VI EPF
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|Brockamp, 1959
Data DOI|
Science Reference|
Science DOI|
Date|1959
Longitude [°E]|-48.2625
Latitude [°N]|69.6981
Location source|Heuberger, 1954
Depth of top measurement [m]|20.0
Depth of bottom measurement [m]|130
Ice thickness [m]|1389
Coverage [% of thickness]|8
Ice thickness source|BedMachine_V3
General_Note|
Temperature_note|Digitized from https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/files/7185520/Polarforsch1965_1-2_8.pdf
Thickness_note|Assuming same location as Heuberger (1954) and CampVI borehole
Location_note|Assuming same location as Heuberger (1954) and CampVI borehole
