Name|penny
Alternate name|Penny Ice Cap
Data source|WIC
Drill year(s)|
Data year(s)|1996
Longitude [°E]|-65.2
Latitude [°N]|67.3
Approximate location name|
Location source|
Ice thickness [m]|176
Ice thickness year|
Ice thickness source|Data file + WIC email (see also Fisher 1998)
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|176.0
