Borehole ID|harrington_2015_46km-11A
Descriptive Name|46km-11A
Area|
Data reference|T. Meierbachtol email
Data DOI|
Science reference|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A948
Date|2011
Longitude [°E]|-49.288804
Latitude [°N]|67.201432
Location source|T. Meierbachtol email
Depth of top measurement [m]|1.0
Depth of bottom measurement [m]|799.0
Ice thickness [m]|821
Coverage [% of thickness]|97
Ice thickness source|T. Meierbachtol email
Measured from: Top, Bottom, Relative|T
General_Note|See data in M1-10 folder
Temperature_note|
Thickness_note|
Location_note|Harrington 2015 name: S5-A
