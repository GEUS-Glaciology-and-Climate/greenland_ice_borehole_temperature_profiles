Borehole ID|grip
Descriptive Name|GRIP
Area|
Data reference|G. Clow email
Data DOI|
Science reference|
Science DOI|
Date|
Longitude [°E]|-37.64
Latitude [°N]|72.58
Location source|Vinther, 2008
Depth of top measurement [m]|40.93
Depth of bottom measurement [m]|3028.57
Ice thickness [m]|3028.57
Coverage [% of thickness]|99
Ice thickness source|Data from Gary Clow
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
