Borehole ID|TD1_88
Place name|Paakitsoq
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Lüthi email
Data DOI|
Science Source|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1988-05-19
Longitude [°E]|-50.13
Latitude [°N]|69.45
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|50.0
Depth of bottom measurement [m]|300
Ice thickness [m]|300
Coverage [% of thickness]|83
Ice thickness source|Unknown PDF: Shallow88II.pdf
Note|
