Borehole ID|Meighen67
Place name|Meighen Ice Cap
Geographic location|Canadian Arctic North
Ice type|Ice cap
Data Source|Graphic in science source
Data DOI|
Science Source|Paterson, W. S. B.: A temperature profile through the Meighen ice cap, Arctic Canada , International Association of Scientific Hydrology 79, 440–449, 1968 
Science DOI|
Date|1965
Longitude [°E]|-99.1
Latitude [°N]|79.9
Location Source|See data source
Depth of top measurement [m]|1.0
Depth of bottom measurement [m]|121
Ice thickness [m]|121
Coverage [% of thickness]|99
Ice thickness source|See data source
Note|Location from Geothermal Database
