Name|td42
Alternate name|
Data source|Unknown PDF: See td1
Drill year(s)|
Data year(s)|1991-08-28
Longitude [°E]|-49.683
Latitude [°N]|69.533
Approximate location name|Paakitsoq
Location source|Unknown PDF: See td1
Ice thickness [m]|>600
Ice thickness year|
Ice thickness source|Unknown PDF: See td1
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|3.0
Depth of bottom measurement [m]|493.0
