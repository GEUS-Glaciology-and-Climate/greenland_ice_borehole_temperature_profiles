Borehole ID|td1
Descriptive Name|
Area|Paakitsoq
Data reference|Unknown PDF: Shallow88II.pdf
Data DOI|
Science reference|
Science DOI|
Date|1988-05-19
Longitude [°E]|-50.13
Latitude [°N]|69.45
Location source|Unknown PDF: Shallow88II.pdf
Depth of top measurement [m]|50.0
Depth of bottom measurement [m]|300.0
Ice thickness [m]|300
Coverage [% of thickness]|83
Ice thickness source|Unknown PDF: Shallow88II.pdf
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
