Borehole ID|CampIII_78b
Place Name|Nunap Kigdlinga
Geographic Location|
Ice Type|
Data Reference|Digitization from published graphic from Stauffer, 1979
Data DOI|
Science Reference|
Science DOI|
Date|1978
Longitude [°E]|-50.0917
Latitude [°N]|69.7176
Location source|M. Lüthi email
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|90.0
Ice thickness [m]|
Coverage [% of thickness]|
Ice thickness source|
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/files/7185440/stauffer_1979.pdf
Thickness_note|
Location_note|
