Borehole ID|hanstausen_hare
Descriptive Name|Hans Tausen Hare
Area|
Data reference|Zekollari, Harry, Huybrechts, Philippe, Noël, Brice, van de Berg, Willem Jan, van den Broeke, Michiel R.: Sensitivity, stability and future evolution of the world’s northernmost ice cap, Hans Tausen Iskappe (Greenland) , The Cryosphere 11(2), Copernicus GmbH, 805–825, 3 2017 
Data DOI|
Science reference|
Science DOI|
Date|
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|288.0
Ice thickness [m]|289
Coverage [% of thickness]|96
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|B
General_Note|
Temperature_note|
Thickness_note|
Location_note|
