Borehole ID|harrington_2015_13km-10
Descriptive Name|13km-10
Area|
Data reference|T. Meierbachtol email
Data DOI|
Science reference|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A941
Date|2010
Longitude [°E]|-50.02945
Latitude [°N]|67.191582
Location source|T. Meierbachtol email
Depth of top measurement [m]|3.5
Depth of bottom measurement [m]|559.0
Ice thickness [m]|
Coverage [% of thickness]|#DIV/0!
Ice thickness source|T. Meierbachtol email
Measured from: Top, Bottom, Relative|T
General_Note|See data in M1-10 folder
Temperature_note|
Thickness_note|
Location_note|Harrington 2015 name: S2
