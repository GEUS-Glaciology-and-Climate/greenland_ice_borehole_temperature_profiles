Borehole ID|agassiz77
Descriptive Name|Agassiz 77 borehole 
Area|Agassiz Ice Cap 
Data reference|W. Colgan email
Data DOI|
Science reference|Clarke, G. K. C., Fisher, D. A., Waddington, E. D.: Wind pumping: A potentially significant heat source in ice sheets , The Physical Basis of Ice Sheet Modelling in Proceedings of the Vancouver Symposium, IAHS , volume 170, 169–180, 1987
Science DOI|
Date|?
Longitude [°E]|-73.1
Latitude [°N]|80.7
Location source|Vinther, 2008
Depth of top measurement [m]|11.0
Depth of bottom measurement [m]|341.0
Ice thickness [m]|340.9
Coverage [% of thickness]|97
Ice thickness source|See data source 
Measured from: Top, Bottom, Relative|T 
General_Note|
Temperature_note|
Thickness_note|Ice thickness from data does not match ice thickness from Vinther (2008)
Location_note|Location approximate
