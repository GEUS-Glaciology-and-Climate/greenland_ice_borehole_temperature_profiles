Borehole ID|site_ii
Descriptive Name|Site II
Area|
Data reference|Hansen, B. L., Landauer, J. K.: Some results of ice cap drill hole measurements, Union Geodesique et Geophysique Internationale. Association Internationale d'Hydrologie Scientifique 47, 313–317, 1958 
Data DOI|
Science reference|
Science DOI|
Date|1958 (late June)
Longitude [°E]|-56.066667
Latitude [°N]|76.983333
Location source|WIC Email
Depth of top measurement [m]|
Depth of bottom measurement [m]|
Ice thickness [m]|1851
Coverage [% of thickness]|0
Ice thickness source|BedMachine
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
