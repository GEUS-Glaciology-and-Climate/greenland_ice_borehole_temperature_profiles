Name|renland
Alternate name|Renland
Data source|BMV
Drill year(s)|1988 (Vinther, 2008)
Data year(s)|1988
Longitude [°E]|-26.768
Latitude [°N]|71.306
Approximate location name|
Location source|Email and Vinther (2008)
Ice thickness [m]|324.4
Ice thickness year|
Ice thickness source|Vinther, B. M., Clausen, H. B., Fisher, D. A., Koerner, R. M., Johnsen, S. J., Andersen, K. K., Dahl-Jensen, D., Rasmussen, S. O., Steffensen, J. P., Svensson, A. M.: Synchronizing ice cores from the Renland and Agassiz ice caps to the Greenland Ice Core Chronology , Journal of Geophysical Research 113(D8), American Geophysical Union (AGU), 4 2008 
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|15.0
Depth of bottom measurement [m]|300.0
