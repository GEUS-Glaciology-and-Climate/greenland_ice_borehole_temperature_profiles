Borehole ID|CampVI
Place Name|Camp VI
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|Digitization from published graphic
Data DOI|
Science Reference|Heuberger, J.-C. 1954. Expéditions Polaires Françaises: Missions Paul-Emil Victor. Glaciologie Groenland Volume 1: Forages sur l'inlandsis. Hermann & Cle, Éditeurs. Paris.
Science DOI|
Date|1950
Longitude [°E]|-48.2625
Latitude [°N]|69.6981
Location source|Heuberger, 1954
Depth of top measurement [m]|4.0
Depth of bottom measurement [m]|125.0
Ice thickness [m]|1389
Coverage [% of thickness]|9
Ice thickness source|BedMachine_V3
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/files/7082104/heuberger_1954.pdf
Thickness_note|
Location_note|
