Borehole ID|Devon72
Place name|Devon Ice Cap
Geographic location|Canadian Arctic North
Ice type|Ice cap
Data Source|Graphic in science source
Data DOI|
Science Source|Paterson, W., R. Koerner, D. Fisher et al. 1977. An oxygen-isotope climatic record from the Devon Island ice cap, Arctic Canada. Nature. 266: 508-511.
Science DOI|10.1038/266508a0
Date|1972
Longitude [°E]|-82.3
Latitude [°N]|75.3
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|213
Ice thickness [m]|300
Coverage [% of thickness]|68
Ice thickness source|See data source
Note|
