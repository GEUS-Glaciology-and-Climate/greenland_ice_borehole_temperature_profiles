Borehole ID|TD3_88
Place name|Paakitsoq
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Lüthi email
Data DOI|
Science Source|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1988-08-18
Longitude [°E]|-50.0
Latitude [°N]|69.48
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|20.0
Depth of bottom measurement [m]|350
Ice thickness [m]|350
Coverage [% of thickness]|94
Ice thickness source|Unknown PDF: See td1. Also Phillips (2010)
Note|
