Name|td51
Alternate name|
Data source|Unknown PDF: See td1 and Lüthi (2015)
Drill year(s)|
Data year(s)|1990-06-09
Longitude [°E]|-49.3
Latitude [°N]|69.566
Approximate location name|Paakitsoq / Swiss Camp
Location source|Unknown PDF: See td1 and Lüthi (2015)
Ice thickness [m]|>600
Ice thickness year|
Ice thickness source|Unknown PDF: See td1 and Lüthi (2015)
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|5.0
Depth of bottom measurement [m]|600.0
