Borehole ID|DYE-3
Place name|DYE-3
Geographic location|South Greenland
Ice type|Ice sheet
Data Source|Graphic in science source
Data DOI|
Science Source|Gundestrup, N. and B. Hansen. 1984. Bore-Hole Survey at Dye 3, South Greenland. Journal of Glaciology. 30: 282–288. 
Science DOI|10.3189/S0022143000006109
Date|1983
Longitude [°E]|-43.8167
Latitude [°N]|65.1833
Location Source|See data source
Depth of top measurement [m]|152.0
Depth of bottom measurement [m]|2030
Ice thickness [m]|2038
Coverage [% of thickness]|92
Ice thickness source|See data source
Velocity [m/yr]|9.7
Note|
