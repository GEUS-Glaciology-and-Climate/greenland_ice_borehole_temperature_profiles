Borehole ID|TD3_88
Place Name|Paakitsoq
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|Unknown PDF: See td1. Also Phillips (2010)
Data DOI|
Science Reference|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1988-08-18
Longitude [°E]|-50.0
Latitude [°N]|69.48
Location source|Colgan, 2021
Depth of top measurement [m]|20.0
Depth of bottom measurement [m]|350.0
Ice thickness [m]|350
Coverage [% of thickness]|94
Ice thickness source|Unknown PDF: See td1. Also Phillips (2010)
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
