Name|jakobshavn_center
Alternate name|
Data source|Iken, A., Echelmeyer, Κ., Harrison, W., Funk, M.: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part I. Measurements of temperature and water level in deep boreholes , Journal of Glaciology 39(131), Cambridge University Press (CUP), 15–25, 1993 
Drill year(s)|
Data year(s)|
Longitude [°E]|
Latitude [°N]|
Approximate location name|
Location source|
Ice thickness [m]|2495
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|12.0
Depth of bottom measurement [m]|2410.0
