Borehole ID|Devon72
Place Name|Devon Ice Cap
Geographic Location|Canadian Arctic North
Ice Type|Ice cap
Data Reference|Paterson, W. S. B., Clarke, G. K. C.: Comparison of theoretical and observed temperature profiles in Devon Island ice cap, Canada , Geophysical Journal International 55(3), Oxford University Press (OUP), 615–632, 12 1978 
Data DOI|
Science Reference|Paterson, W., R. Koerner, D. Fisher et al. 1977. An oxygen-isotope climatic record from the Devon Island ice cap, Arctic Canada. Nature. 266: 508-511.
Science DOI|10.1038/266508a0
Date|1972
Longitude [°E]|-82.3
Latitude [°N]|75.3
Location source|Colgan, 2021
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|213.0
Ice thickness [m]|300
Coverage [% of thickness]|68
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
