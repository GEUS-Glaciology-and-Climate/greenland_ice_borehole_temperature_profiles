Borehole ID|ngrip
Descriptive Name|NGRIP
Area|
Data reference|G. Clow email
Data DOI|
Science reference|
Science DOI|
Date|2003
Longitude [°E]|-42.32
Latitude [°N]|75.1
Location source|Vinther (2008)
Depth of top measurement [m]|81.89
Depth of bottom measurement [m]|2992.47
Ice thickness [m]|3085
Coverage [% of thickness]|94
Ice thickness source|See data source email
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
