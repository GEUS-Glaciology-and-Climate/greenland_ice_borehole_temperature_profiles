Borehole ID|Isunnguata_46km-11A
Place name|Isunnguata Sermia
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Meierbachtol email
Data DOI|
Science Source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A948
Date|2011
Longitude [°E]|-49.2888
Latitude [°N]|67.20143
Location Source|Meierbachtol email
Depth of top measurement [m]|1.0
Depth of bottom measurement [m]|799
Ice thickness [m]|821
Coverage [% of thickness]|97
Ice thickness source|T. Meierbachtol email
Note|See data in M1-10 folder; Harrington 2015 name: S5-A
