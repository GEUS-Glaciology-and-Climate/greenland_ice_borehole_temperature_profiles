Name|td7
Alternate name|
Data source|Tech Report
Drill year(s)|
Data year(s)|
Longitude [°E]|
Latitude [°N]|
Approximate location name|
Location source|
Ice thickness [m]|
Ice thickness year|
Ice thickness source|
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|
Depth of bottom measurement [m]|
