Borehole ID|Devon98
Place Name|Devon Ice Cap
Geographic Location|Canadian Arctic North
Ice Type|Cap
Data Reference|W. Colgan email
Data DOI|
Science Reference|Paterson, W., R. Koerner, D. Fisher et al. 1977. An oxygen-isotope climatic record from the Devon Island ice cap, Arctic Canada. Nature. 266: 508-511.
Science DOI|10.1038/266508a0
Date|2000-04-15
Longitude [°E]|-82.3
Latitude [°N]|75.3
Location source|Colgan2021
Depth of top measurement [m]|13.0
Depth of bottom measurement [m]|218.0
Ice thickness [m]|301.0
Coverage [% of thickness]|68
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
