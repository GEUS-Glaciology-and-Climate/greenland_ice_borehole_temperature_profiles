Borehole ID|Devon98
Place name|Devon Ice Cap
Geographic location|Canadian Arctic North
Site type|Ice cap
Data Source|Zdanowicz email
Data DOI|
Science Source|Kinnard, C., C. Zdanowicz, D. Fisher et al. 2006. Calibration of an ice-core glaciochemical (sea-salt) record with Sea-ice variability in the Canadian Arctic. Annals of Glaciology. 44: 383-390. 
Science DOI|10.3189/172756406781811349
Date|2000-04-15
Longitude [°E]|-82.3
Latitude [°N]|75.3
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|13.0
Depth of bottom measurement [m]|218
Ice thickness [m]|301
Coverage [% of thickness]|68
Ice thickness source|See data source
Note|
