Name|h2015_s1b
Alternate name|
Data source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Drill year(s)|
Data year(s)|2011-2013
Longitude [°E]|
Latitude [°N]|
Approximate location name|
Location source|
Ice thickness [m]|145
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|6.0
Depth of bottom measurement [m]|131.0
