Borehole ID|SiteII
Place name|Site II
Geographic location|Northwest Greenland
Site type|Ice sheet
Data Source|Graphic in science source
Data DOI|
Science Source|Hansen, B. and J. Landauer. 1958. Some results of ice cap drill hole measurements. IASH Publication. 47: 313-317.
Science DOI|
Date|1958-06-25
Longitude [°E]|-56.07
Latitude [°N]|76.98
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|16.0
Depth of bottom measurement [m]|410
Ice thickness [m]|1851
Coverage [% of thickness]|21
Ice thickness source|BedMachine_V3
Note|
