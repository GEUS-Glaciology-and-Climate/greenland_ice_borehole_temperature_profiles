Borehole ID|devon_72
Descriptive Name|Devon borehole
Area|Devon Ice Cap
Data reference|Paterson, W. S. B., Clarke, G. K. C.: Comparison of theoretical and observed temperature profiles in Devon Island ice cap, Canada , Geophysical Journal International 55(3), Oxford University Press (OUP), 615–632, 12 1978 
Data DOI|
Science reference|
Science DOI|
Date|
Longitude [°E]|-82.14
Latitude [°N]|75.34
Location source|
Depth of top measurement [m]|9.0
Depth of bottom measurement [m]|299.0
Ice thickness [m]|299
Coverage [% of thickness]|97
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
