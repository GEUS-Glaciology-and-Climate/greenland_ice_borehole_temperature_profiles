Borehole ID|GISP2
Place name|GISP2
Geographic location|Central Greenland
Ice type|Ice sheet
Data Source|Clow email
Data DOI|
Science Source|MacGregor, J., J. Li, J. Paden et al. 2015. Radar attenuation and temperature within the Greenland Ice Sheet. Journal of Geophysical Research. 120: 983-1008. 
Science DOI|10.1002/2014JF003418
Date|1996-06-02
Longitude [°E]|-38.4667
Latitude [°N]|72.5833
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|73.0
Depth of bottom measurement [m]|3053
Ice thickness [m]|3053
Coverage [% of thickness]|98
Ice thickness source|https://en.wikipedia.org/wiki/List_of_ice_cores#Greenland
Velocity [m/yr]|1.7
Note|Ice thickness from data does not match ice thickness from Vinther (2008); Location approximate
