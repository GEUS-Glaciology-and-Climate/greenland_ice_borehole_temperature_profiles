Name|camp_vi
Alternate name|Camp VI
Data source|Lüthi pers. comm -> Heuberger (1950) p. 47, 31.1
Drill year(s)|1950?
Data year(s)|1950?
Longitude [°E]|
Latitude [°N]|
Approximate location name|
Location source|
Ice thickness [m]|
Ice thickness year|
Ice thickness source|
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|4
Depth of bottom measurement [m]|125
