Borehole ID|td51
Descriptive Name|
Area|Paakitsoq / Swiss Camp
Data reference|Unknown PDF: See td1 and Lüthi (2015)
Data DOI|
Science reference|
Science DOI|
Date|1990-06-09
Longitude [°E]|-49.3
Latitude [°N]|69.566
Location source|Unknown PDF: See td1 and Lüthi (2015)
Depth of top measurement [m]|5.0
Depth of bottom measurement [m]|600.0
Ice thickness [m]|>600
Coverage [% of thickness]|#VALUE!
Ice thickness source|Unknown PDF: See td1 and Lüthi (2015)
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
