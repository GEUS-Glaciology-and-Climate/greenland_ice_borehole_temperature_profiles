Borehole ID|Barnes_T020_1979
Place name|Barnes Ice Cap
Geographic location|Canadian Arctic South
Ice type|Ice cap
Data Source|Graphic in science source
Data DOI|
Science Source|Hooke, Roger LeB., Alexander, E. Calvin, Gustafson, Robert J.: Temperature profiles in the Barnes Ice Cap, Baffin Island, Canada, and heat flux from the subglacial terrane , Canadian Journal of Earth Sciences 17(9), Canadian Science Publishing, 1174–1188, sep 1980
Science DOI|10.1139/e80-124
Date|1979-07-02
Longitude [°E]|-71.892
Latitude [°N]|69.71965
Location Source|Location digitized by M. Jacquemart from Gilbert (2016) and Hooke (1980)
Depth of top measurement [m]|0.0
Depth of bottom measurement [m]|279
Ice thickness [m]|369
Coverage [% of thickness]|76
Ice thickness source|Hooke, Roger LeB., Alexander, E. Calvin, Gustafson, Robert J.: Temperature profiles in the Barnes Ice Cap, Baffin Island, Canada, and heat flux from the subglacial terrane , Canadian Journal of Earth Sciences 17(9), Canadian Science Publishing, 1174–1188, sep 1980
Note|"Date is ""Date completed"" from Hooke (1980) Table 1 Column 2 + Days to final measurement (Column 3); Location digitized by M. Jacquemart"
