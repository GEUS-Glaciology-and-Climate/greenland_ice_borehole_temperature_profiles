Borehole ID|Barnes_14.3_T_1975
Place name|Barnes Ice Cap
Geographic location|Canadian Arctic South
Ice type|Ice cap
Data Source|Table in science source
Data DOI|
Science Source|Classen, D. F.: Temperature profiles for the Barnes Ice Cap surge zone , Journal of Glaciology 18(80), International Glaciological Society, 391–405, 1977
Science DOI|10.3189/s0022143000021079
Date|1975-07-02
Longitude [°E]|-72.1495
Latitude [°N]|69.63971832
Location Source|See Science Source
Depth of top measurement [m]|140.0
Depth of bottom measurement [m]|200
Ice thickness [m]|220
Coverage [% of thickness]|27
Ice thickness source|See science source
Note|Location digitized by M. Jacquemart
