Site|Alternate name|Data source|Data year(s)|Depth of top measurement [m]|Depth of bottom measurement [m]|Drill year(s)|Longitude [°E]|Latitude [°N]|Approximate location name|Location source|Ice thickness [m]|Ice thickness year|Ice thickness source|Surface velocity [m yr^-1]|Surface velocity year|Surface velocity source|Measured from: Top, Bottom, Relative|Coverage [% of thickness]
agassiz77|Agassiz 77 borehole |WIC Email|1977|11.0 |341.0 |1977 (Vinther, 2008)|-73.1 |80.7 |Agassiz Ice Cap |Vinther, 2008|340.9 ||See data source ||||T |97
agassiz79a|Agassiz ice cap 1979A borehole |WIC Email |1979 |12.0 |142.0 |1979 (Vinther, 2008)|-73.1 |80.7 |Agassiz Ice Cap |Vinther, 2008|141.9 |nan |See data source |nan |nan |nan |T |92
agassiz79b|Agassiz ice cap 1979B borehole|WIC Email|1979|11.0|141.0|1979 (Vinther, 2008)|-73.1|80.7|Agassiz Ice Cap|Vinther (2008)|141.2||See data source||||T|92
agassiz84|Agassiz 1984 borehole|WIC Email|1984|3.0|128.0|184 (Vinther, 2008)|-73.1|80.7|Agassiz Ice Cap|Vinther, 2008|127.6||See data source||||T|98
camp_century|Camp Century|Weertman, J.: Comparison betwe||9.0|1387.0||||Camp Century|?|1387|?|?||||B|99
camp_vi|Camp VI|Lüthi pers. comm -> Heuberger (1950) p. 47, 31.1|1950?|4|125|1950?|||||||||||T|0
devon_00|Devon borehole|WIC Email|2000-04-15|13|218|1998-04-15 to 1998-05-07|-82.14|75.34|Devon Ice Cap||300.55||See data source||||T|68
devon_71|Devon borehole|Paterson, W. S. B., Clarke, G. K. C.: Comparison of theoretical and observed temperature profiles in Devon Island ice cap, Canada , Geophysical Journal International 55(3), Oxford University Press (OUP), 615–632, 12 1978 ||10|213||||Devon Ice Cap||300|drill year|See data source||||T|68
devon_72|Devon borehole|Paterson, W. S. B., Clarke, G. K. C.: Comparison of theoretical and observed temperature profiles in Devon Island ice cap, Canada , Geophysical Journal International 55(3), Oxford University Press (OUP), 615–632, 12 1978 ||9|299||-82.14|75.34|Devon Ice Cap||299|drill year|See data source||||T|97
dye_3|DYE-3|Gundestrup, N. S., Hansen, B. Lyle: Bore-Hole Survey at Dye 3, South Greenland , Journal of Glaciology 30(106), Cambridge University Press (CUP), 282–288, 1984 |1983|152|2030|1979 to 1981|-43.816667|65.183333|South Greenland|See data source|2038|1983|See data source||||T|92
flade_isblink|Flade Isblink|Dorthe Dalh-Jensen (personal comm.)||80.0|420.0||-15.7029|81.2926|||540||See WIC email||||T|63
foxx1|FOXX|Lüthi, Martin P., Ryser, Claudia, Andrews, Lauren C., Catania, Ginny A., Funk, Martin, Hawley, Robert L., Hoffman, Matthew J., Neumann, Thomas A.: Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming , The Cryosphere 9(1), 245–253, 2015 |2011-2013|6|611||||Paakitsoq||631||See data source||||T|96
foxx2|FOXX2|Lüthi, Martin P., Ryser, Claudia, Andrews, Lauren C., Catania, Ginny A., Funk, Martin, Hawley, Robert L., Hoffman, Matthew J., Neumann, Thomas A.: Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming , The Cryosphere 9(1), 245–253, 2015 |2011-2013|8.6|285.9||||Paakitsoq||||||||T|0
gisp2|GISP2; GISP II|Cuffey, Kurt M., Alley, Richard B., Grootes, Pieter M., Anandakrishnan, Sridhar: Toward using borehole temperatures to calibrate an isotopic paleothermometer in central Greenland , Palaeogeography, Palaeoclimatology, Palaeoecology 98(2-4), Elsevier BV, 265–268, 12 1992 |1989,1990|37.0|216.0||||Russell / Leverett ?||3100||Hodge 1990?||||T|6
grip|GRIP|Johnsen, Sigfus J., Dahl-Jensen, Dorthe, Dansgaard, Willi, Gundestrup, Niels: Greenland palaeotemperatures derived from GRIP bore hole temperature and ice core isotope profiles , Tellus B: Chemical and Physical Meteorology 47(5), Informa UK Limited, 624–629, 1 1995 ||107.0|3023.0|1989-1992 (Vinther, 2008)|-37.64|72.58||Vinther (2008)|3027||Montagnat, M., Azuma, N., Dahl-Jensen, D., Eichler, J., Fujita, S., Gillet-Chaulet, F., Kipfstuhl, S., Samyn, D., Svensson, A., Weikusat, I.: Fabric along the NEEM ice core, Greenland, and its comparison with GRIP and NGRIP ice cores , The Cryosphere 8(4), Copernicus GmbH, 1129–1138, 7 2014 ||||T|96
gull|GULL|Lüthi, Martin P., Ryser, Claudia, Andrews, Lauren C., Catania, Ginny A., Funk, Martin, Hawley, Robert L., Hoffman, Matthew J., Neumann, Thomas A.: Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming , The Cryosphere 9(1), 245–253, 2015 |2011-2013|4|704||||Paakitsoq||703||See data source||||T|100
h2015_s1a||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|11.0|81.0||||||92||See data source||||T|76
h2015_s1b||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|6.0|131.0||||||145||See data source||||T|86
h2015_s2a||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|3.5|559||||||||See data source||||T|0
h2015_s3a||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|218.0|368.0||||||458||See data source||||T|33
h2015_s3b||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|27.0|460.0||||||466||See data source||||T|93
h2015_s3c||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|20.0|459.0||||||460||See data source||||T|95
h2015_s4a||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|11.0|690.0||||||701||See data source||||T|97
h2015_s4b||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|18.0|690.0||||||692||See data source||||T|97
h2015_s4c||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|17.0|688.0||||||698||See data source||||T|96
h2015_s5a||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|1.0|799.0||||||821||See data source||||T|97
h2015_s5b||Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 |2011-2013|114.0|728.0||||||815||See data source||||T|75
hanstausen_dome|Hans Tausen Dome|Zekollari, Harry, Huybrechts, Philippe, Noël, Brice, van de Berg, Willem Jan, van den Broeke, Michiel R.: Sensitivity, stability and future evolution of the world’s northernmost ice cap, Hans Tausen Iskappe (Greenland) , The Cryosphere 11(2), Copernicus GmbH, 805–825, 3 2017 ||10.0|344.0||||||345||See data source||||B|97
hanstausen_hare|Hans Tausen Hare|Zekollari, Harry, Huybrechts, Philippe, Noël, Brice, van de Berg, Willem Jan, van den Broeke, Michiel R.: Sensitivity, stability and future evolution of the world’s northernmost ice cap, Hans Tausen Iskappe (Greenland) , The Cryosphere 11(2), Copernicus GmbH, 805–825, 3 2017 ||10.0|288.0||||||289||See data source||||B|96
isua_10|Isua|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 |1972-1973|5.0|95.0||-49.75|65.2093|||97||See data source||||T|93
isua_11|Isua|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 |1972-1973|25.0|116.0||-49.7510|65.2072|||120||See data source||||T|76
isua_12|Isua|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 |1972-1973|25.0|95.0||-49.753|65.2039|||100||See data source||||T|70
isua_13|Isua|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 |1972-1973|6.0|247.0||-49.7456|65.2069|||265||See data source||||T|91
isua_14|Isua|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 |1972-1973|6.0|237.0||-49.7443|65.2058|||299||See data source||||T|77
jakobshavn_center||Iken, A., Echelmeyer, Κ., Harrison, W., Funk, M.: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part I. Measurements of temperature and water level in deep boreholes , Journal of Glaciology 39(131), Cambridge University Press (CUP), 15–25, 1993 ||12.0|2410.0||||||2495||See data source||||T|96
jakobshavn_left||Iken, A., Echelmeyer, Κ., Harrison, W., Funk, M.: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part I. Measurements of temperature and water level in deep boreholes , Journal of Glaciology 39(131), Cambridge University Press (CUP), 15–25, 1993 ||8.0|1517.0||||||1530||See data source||||T|99
jakobshavn_sheet||Lüthi, Martin, Funk, Martin, Iken, Almut, Gogineni, Shivaprasad, Truffer, Martin: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part III. Measurements of ice deformation, temperature and cross-borehole conductivity in boreholes to the bedrock , Journal of Glaciology 48(162), 369–385, 2002 ||19.0|798.0||||||828||See data source||||T|94
m2020_14n||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|37.0|647.0||||||660||See data source||||B|92
m2020_14sa||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|58.0|659.0||||||660||See data source||||B|91
m2020_14sb||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|499.0|650.0||||||660||See data source||||B|23
m2020_14w||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|39.0|659.0||||||660||See data source||||B|94
m2020_15ca||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|35.0|654.0||||||660||See data source||||B|94
m2020_15cb||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|355.0|655.0||||||660||See data source||||B|45
m2020_15e||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|35.0|656.0||||||660||See data source||||B|94
m2020_15n||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|35.0|655.0||||||660||See data source||||B|94
m2020_15s||McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 |2017|35.0|655.0||||||660||See data source||||B|94
meighan|Meighan Ice Cap|Paterson, W. S. B.: A temperature profile through the Meighen ice cap, Arctic Canada , International Association of Scientific Hydrology 79, 440–449, 1968 |1965|1.0|121.0||||||121.2||See data source||||T|99
neem|NEEM|MacGregor, Joseph A., Li, Jilu, Paden, John D., Catania, Ginny A., Clow, Gary D., Fahnestock, Mark A., Gogineni, S. Prasad, Grimm, Robert E., Morlighem, Mathieu, Nandi, Soumyaroop, et al.: Radar attenuation and temperature within the Greenland Ice Sheet , Journal of Geophysical Research: Earth Surface 120(6), American Geophysical Union (AGU), 983–1008, 6 2015 ||91.0|2509.0|2008 through 2012|-51.06|77.45|Northwest Greenland|Dahl-Jensen, D., Albert, Mary R., Aldahan, A., Azuma, N., Balslev-Clausen, D., Baumgartner, M., Berggren, A. -M., Bigler, M., Binder, T., Blunier, T., Bourgeois, J. C., Brook, E. J., Buchardt, S. L., Buizert, C., Capron, E., Chappellaz, J., Chung, J., Clausen, H. B., Cvijanovic, I., Davies, S. M., Ditlevsen, P., Eicher, O., Fischer, H., Fisher, D. A., Fleet, L. G., Gfeller, G., Gkinis, V., Gogineni, S., Goto-Azuma, K., Grinsted, A., Gudlaugsdottir, H., Guillevic, M., Hansen, S. B., Hansson, M., Hirabayashi, M., Hong, S., Hur, S. D., Huybrechts, Philippe, Hvidberg, C. S., Iizuka, Y., Jenk, T., Johnsen, S. J., Jones, T. R., Jouzel, J., Karlsson, N. B., Kawamura, K., Keegan, K., Kettner, E., Kipfstuhl, S., Kjær, H. A., Koutnik, M., Kuramoto, T., Koehler, P., Laepple, T., Landais, A., Langen, P. L., Larsen, L. B., Leuenberger, D., Leuenberger, M., Leuschen, C., Li, J., Lipenkov, V., Martinerie, P., Maselli, O. J., Masson-Delmotte, V., McConnell, J. R., Miller, H., Mini, O., Miyamoto, A., Montagnat-Rentier, M., Mulvaney, R., Muscheler, Raimund, Orsi, A. J., Paden, J., Panton, C., Pattyn, F., Petit, J. -R., Pol, K., Popp, T., Possnert, G., Prie, F., Prokopiou, M., Quiquet, A., Rasmussen, S. O., Raynaud, D., Ren, J., Reutenauer, C., Ritz, C., Rockmann, T., Rosen, J. L., Rubino, M., Rybak, O., Samyn, D., Sapart, C. J., Schilt, A., Schmidt, A. M. Z., Schwander, J., Schuepbach, S., Seierstad, I., Severinghaus, J. P., Sheldon, S., Simonsen, S. B., Sjolte, Jesper, Solgaard, A. M., Sowers, T., Sperlich, P., Steen-Larsen, H. C., Steffen, K., Steffensen, J. P., Steinhage, D., Stocker, T. F., Stowasser, C., Sturevik, A. S., Sturges, W. T., Sveinbjornsdottir, A., Svensson, A., Tison, J. -L., Uetake, J., Vallelonga, P., van de Wal, R. S. W., van der Wel, G., Vaughn, B. H., Vinther, B., Waddington, E., Wegner, A., Weikusat, I., White, J. W. C., Wilhelms, F., Winstrup, M., Witrant, E., Wolff, E. W., Xiao, C., Zheng, J.: Eemian interglacial reconstructed from a Greenland folded ice core , Nature 493(7433), Nature Publishing Group, 489–494, 2013 |2538||MacGregor, Joseph A., Fahnestock, Mark A., Catania, Ginny A., Aschwanden, Andy, Clow, Gary D., Colgan, William T., Gogineni, Prasad S., Morlighem, Mathieu, Nowicki, Sophie M. J., Paden, John D., Price, Stephen F., Seroussi, Hélène: A synthesis of the basal thermal state of the Greenland Ice Sheet , Journal of Geophysical Research: Earth Surface 121(7), 1328–1350, 2016 ||||R|95
ngrip|NGRIP|Dahl-Jensen, Dorthe, Gundestrup, Niels, Gogineni, S Prasad, Miller, Heinz: Basal melt at NorthGRIP modeled from borehole, ice-core and radio-echo sounder observations , Annals of Glaciology 37, International Glaciological Society, 207–212, 2003 ||204.0|2888.0|1996-2004 (Vinther, 2008)|-42.32|75.10||Vinther (2008)|3080||See data source||||T|87
penny|Penny Ice Cap|WIC|1996|10.0|176.0||-65.2|67.3|||176||Data file + WIC email (see also Fisher 1998)||||T|94
pow|Prince of Wales|WIC|2005-05-15|10.0|176.0||-80.395|78.3897|||176||WIC||||T|94
renland|Renland|BMV|1988|15.0|300.0|1988 (Vinther, 2008)|-26.768|71.306||Email and Vinther (2008)|324.4||Vinther, B. M., Clausen, H. B., Fisher, D. A., Koerner, R. M., Johnsen, S. J., Andersen, K. K., Dahl-Jensen, D., Rasmussen, S. O., Steffensen, J. P., Svensson, A. M.: Synchronizing ice cores from the Renland and Agassiz ice caps to the Greenland Ice Core Chronology , Journal of Geophysical Research 113(D8), American Geophysical Union (AGU), 4 2008 ||||T|88
site_ii|Site II|Hansen, B. L., Landauer, J. K.: Some results of ice cap drill hole measurements, Union Geodesique et Geophysique Internationale. Association Internationale d'Hydrologie Scientifique 47, 313–317, 1958 |1958 (late June)|||1957 (Summer)|-56.066667|76.983333||WIC Email|1851||BedMachine||||T|0
td1||Unknown PDF: Shallow88II.pdf|1988-05-19|50.0|300.0||-50.13|69.45|Paakitsoq|Unknown PDF: Shallow88II.pdf|300||Unknown PDF: Shallow88II.pdf||||T|83
td2||Unknown PDF: See td1|1988-05-19|27.0|202.0||-50.13|69.45|Paakitsoq|Unknown PDF: See td1|470||Unknown PDF: See td1||||T|37
td3||Unknown PDF: See td1. Also Phillips (2010)|1988-08-18|20.0|350.0||-50.00|69.483|Paakitsoq|Unknown PDF: See td1. Also Phillips (2010)|350||Unknown PDF: See td1. Also Phillips (2010)||||T|94
td41||Unknown PDF: See td1|1991-11-05|5.0|495.0||-49.683|69.533|Paakitsoq|Unknown PDF: See td1|>600||Unknown PDF: See td1||||T|0
td42||Unknown PDF: See td1|1991-08-28|3.0|493.0||-49.683|69.533|Paakitsoq|Unknown PDF: See td1|>600||Unknown PDF: See td1||||T|0
td51||Unknown PDF: See td1 and Lüthi (2015)|1990-06-09|5.0|600.0||-49.3|69.566|Paakitsoq / Swiss Camp|Unknown PDF: See td1 and Lüthi (2015)|>600||Unknown PDF: See td1 and Lüthi (2015)||||T|0
td52||Unknown PDF: See td1 and Lüthi (2015)|1991-05-25|5.0|600.0||-49.3|69.566|Paakitsoq / Swiss Camp|Unknown PDF: See td1 and Lüthi (2015)|>600||Unknown PDF: See td1 and Lüthi (2015)||||T|0
td6||Tech Report|||||||||||||||T|0
td7||Tech Report|||||||||||||||T|0
td8||Tech Report|||||||||||||||T|0
tuto_ramp|Tuto Ramp|Davis, RM: Approach roads, Greenland 1960–1964 , Technical Report 133. Corps of Engineers, Cold Regions Research & Engineering Laboratory , 1967 |1962 (August)||||-68.287295|76.41133|Thule Approach Road(?)||48||See data source|1.0||WIC Email|T(ish)|0
