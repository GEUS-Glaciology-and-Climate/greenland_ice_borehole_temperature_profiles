Name|pow
Alternate name|Prince of Wales
Data source|WIC
Drill year(s)|
Data year(s)|2005-05-15
Longitude [°E]|-80.395
Latitude [°N]|78.3897
Approximate location name|
Location source|
Ice thickness [m]|176
Ice thickness year|
Ice thickness source|WIC
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|176.0
