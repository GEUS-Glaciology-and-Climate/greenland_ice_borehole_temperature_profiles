Borehole ID|PrinceWales05
Place Name|Prince of Wales Ice Cap
Geographic Location|Canadian Arctic North
Ice Type|
Data Reference|W. Colgan email
Data DOI|
Science Reference|Kinnard, C., R. Koerner, C. Zdanowicz et al. 2008. Stratigraphic analysis of an ice core from the Prince of Wales Icefield, Ellesmere Island, Arctic Canada, using digital image analysis: High‐resolution density, past summer warmth reconstruction, and melt effect on ice core solid conductivity. Journal of Geophysical Research. 113: D24120. 
Science DOI|10.1029/2008JD011083
Date|2005-05-15
Longitude [°E]|-80.395
Latitude [°N]|78.3897
Location source|Colgan2021
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|176.0
Ice thickness [m]|176.0
Coverage [% of thickness]|94
Ice thickness source|WIC
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
