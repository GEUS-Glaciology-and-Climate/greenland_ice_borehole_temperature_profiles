Borehole ID|hills_2017_15n
Descriptive Name|33km_15N
Area|Isunnguata Sermia
Data reference|Joel Harper. 2017. Ice temperatures measured in a grid of boreholes, Western Greenland, 2014-2016. Arctic Data Center. doi:10.18739/A24746S04.
Data DOI|10.18739/A24746S04
Science reference|"Hills, Benjamin H., Joel T. Harper, Neil F. Humphrey, and Toby W. Meierbachtol. ""Measured horizontal temperature gradients constrain heat transfer mechanisms in Greenland ice."" Geophysical Research Letters 44, no. 19 (2017): 9778-9785."
Science DOI|10.1002/2017GL074917
Date|2016
Longitude [°E]|-49.566914
Latitude [°N]|67.18312399999999
Location source|10.18739/A24746S04
Depth of top measurement [m]|15.0
Depth of bottom measurement [m]|635.0
Ice thickness [m]|640
Coverage [% of thickness]|97
Ice thickness source|10.18739/A24746S04
Measured from: Top, Bottom, Relative|B
General_Note|See also McDowell, I. E., Humphrey, N. F., Harper, J. T., and Meierbachtol, T. W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet, The Cryosphere, 15, 897–907, https://doi.org/10.5194/tc-15-897-2021, 2021.
Temperature_note|
Thickness_note|
Location_note|
