Name|td2
Alternate name|
Data source|Unknown PDF: See td1
Drill year(s)|
Data year(s)|1988-05-19
Longitude [°E]|-50.13
Latitude [°N]|69.45
Approximate location name|Paakitsoq
Location source|Unknown PDF: See td1
Ice thickness [m]|470
Ice thickness year|
Ice thickness source|Unknown PDF: See td1
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|27.0
Depth of bottom measurement [m]|202.0
