Borehole ID|CampVI_50
Place name|Camp VI
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Table in science source
Data DOI|
Science Source|Heuberger, J.-C. 1954. Expéditions Polaires Françaises: Missions Paul-Emil Victor. Glaciologie Groenland Volume 1: Forages sur l'inlandsis. Hermann & Cle, Éditeurs. Paris.
Science DOI|
Date|1950
Longitude [°E]|-48.2625
Latitude [°N]|69.6981
Location Source|Heuberger, 1954
Depth of top measurement [m]|4.0
Depth of bottom measurement [m]|125
Ice thickness [m]|1389
Coverage [% of thickness]|9
Ice thickness source|BedMachine_V3
Velocity [m/yr]|154.8
Note|
