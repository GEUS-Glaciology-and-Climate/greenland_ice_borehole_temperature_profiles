Borehole ID|HansTausen_Hare
Place name|Hans Tausen Hare
Geographic location|North Greenland
Ice type|Ice cap
Data Source|Zekollari email
Data DOI|
Science Source|Zekollari, Harry, Huybrechts, Philippe, Noël, Brice, van de Berg, Willem Jan, van den Broeke, Michiel R.: Sensitivity, stability and future evolution of the world’s northernmost ice cap, Hans Tausen Iskappe (Greenland) , The Cryosphere 11(2), Copernicus GmbH, 805–825, 3 2017 
Science DOI|10.5194/tc-11-805-2017
Date|1995
Longitude [°E]|-36.67
Latitude [°N]|82.84
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|9.0
Depth of bottom measurement [m]|288
Ice thickness [m]|289
Coverage [% of thickness]|97
Ice thickness source|See data source
Note|Drill date: 10.34194/bullggu.v172.6749 
