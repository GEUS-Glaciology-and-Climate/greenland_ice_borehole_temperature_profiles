Name|td3
Alternate name|
Data source|Unknown PDF: See td1. Also Phillips (2010)
Drill year(s)|
Data year(s)|1988-08-18
Longitude [°E]|-50.00
Latitude [°N]|69.483
Approximate location name|Paakitsoq
Location source|Unknown PDF: See td1. Also Phillips (2010)
Ice thickness [m]|350
Ice thickness year|
Ice thickness source|Unknown PDF: See td1. Also Phillips (2010)
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|20.0
Depth of bottom measurement [m]|350.0
