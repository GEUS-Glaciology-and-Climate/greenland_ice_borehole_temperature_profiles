Borehole ID|flade_isblink
Descriptive Name|Flade Isblink
Area|
Data reference|Dorthe Dalh-Jensen (personal comm.)
Data DOI|
Science reference|
Science DOI|
Date|
Longitude [°E]|-15.7029
Latitude [°N]|81.2926
Location source|
Depth of top measurement [m]|80.0
Depth of bottom measurement [m]|420.0
Ice thickness [m]|540
Coverage [% of thickness]|63
Ice thickness source|See WIC email
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
