Borehole ID|DYE-3
Place Name|DYE-3
Geographic Location|South Greenland
Ice Type|Ice sheet
Data Reference|Gundestrup, N. S., Hansen, B. Lyle: Bore-Hole Survey at Dye 3, South Greenland , Journal of Glaciology 30(106), Cambridge University Press (CUP), 282–288, 1984 
Data DOI|
Science Reference|Gundestrup, N. and B. Hansen. 1984. Bore-Hole Survey at Dye 3, South Greenland. Journal of Glaciology. 30: 282–288. 
Science DOI|10.3189/S0022143000006109
Date|1983
Longitude [°E]|-43.8167
Latitude [°N]|65.1833
Location source|See data source
Depth of top measurement [m]|152.0
Depth of bottom measurement [m]|2030
Ice thickness [m]|2038
Coverage [% of thickness]|92
Ice thickness source|See data source
General_Note|
Temperature_note|
Thickness_note|
Location_note|
