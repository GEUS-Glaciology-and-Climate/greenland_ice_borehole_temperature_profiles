Borehole ID|Jakobshavn95D_I1
Place name|Jakobshavn Isbræ
Geographic location|Central West Greenland
Site type|Ice sheet
Data Source|Lüthi email
Data DOI|
Science Source|Lüthi, Martin, Funk, Martin, Iken, Almut, Gogineni, Shivaprasad, Truffer, Martin: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part III. Measurements of ice deformation, temperature and cross-borehole conductivity in boreholes to the bedrock, Journal of Glaciology 48(162), 369–385, 2002 
Science DOI|10.3189/172756502781831322
Date|1995
Longitude [°E]|-48.6869
Latitude [°N]|69.235
Location Source|10.3189/172756502781831322
Depth of top measurement [m]|344.0
Depth of bottom measurement [m]|829
Ice thickness [m]|832
Coverage [% of thickness]|58
Ice thickness source|See science reference
Note|
