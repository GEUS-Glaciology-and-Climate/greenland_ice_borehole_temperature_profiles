Borehole ID|Isunnguata_27km-12C
Place name|Isunnguata Sermia
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Meierbachtol email
Data DOI|
Science Source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A947
Date|2012
Longitude [°E]|-49.71811
Latitude [°N]|67.20382
Location Source|T. Meierbachtol email
Depth of top measurement [m]|17.0
Depth of bottom measurement [m]|688
Ice thickness [m]|696
Coverage [% of thickness]|96
Ice thickness source|T. Meierbachtol email
Note|See data in M1-10 folder; Harrington 2015 name: S4-C
