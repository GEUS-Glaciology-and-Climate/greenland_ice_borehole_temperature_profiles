Borehole ID|TD4_91a
Place Name|Paakitsoq
Geographic Location|Central West Greenland
Ice Type|
Data Reference|Unknown PDF: See td1
Data DOI|
Science Reference|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1991-11-05
Longitude [°E]|-49.68
Latitude [°N]|69.53
Location source|Colgan2021
Depth of top measurement [m]|5.0
Depth of bottom measurement [m]|495.0
Ice thickness [m]|600.0
Coverage [% of thickness]|82
Ice thickness source|Estimate. lower bound Unknown PDF, upper bound BedMachine_V3
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
