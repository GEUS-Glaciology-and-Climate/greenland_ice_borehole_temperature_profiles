Borehole ID|Jakobshavn89B
Place Name|Jakobshavn Isbræ
Geographic Location|Central West Greenland
Ice Type|
Data Reference|M. Lüthi email
Data DOI|
Science Reference|Iken, A., Echelmeyer, Κ., Harrison, W., Funk, M.: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part I. Measurements of temperature and water level in deep boreholes , Journal of Glaciology 39(131), Cambridge University Press (CUP), 15–25, 1993 
Science DOI|10.3189/S0022143000015689
Date|1989
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|
Depth of bottom measurement [m]|
Ice thickness [m]|2520.0
Coverage [% of thickness]|100
Ice thickness source|See science reference
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
