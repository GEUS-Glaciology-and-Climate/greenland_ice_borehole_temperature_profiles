Borehole ID|Isunnguata_M1-10
Place name|Isunnguata Sermia
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Meierbachtol email
Data DOI|
Science Source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A939
Date|2010
Longitude [°E]|-50.06427
Latitude [°N]|67.16221
Location Source|T. Meierbachtol email
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|90
Ice thickness [m]|99
Coverage [% of thickness]|81
Ice thickness source|T. Meierbachtol email
Note|See data in M1-10 folder; Harrington 2015 name: S1-A
