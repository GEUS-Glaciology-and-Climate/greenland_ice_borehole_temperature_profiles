Borehole ID|h2015_s4b
Descriptive Name|27km_S4B
Area|
Data reference|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Data DOI|
Science reference|
Science DOI|
Date|2012
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|18.0
Depth of bottom measurement [m]|690.0
Ice thickness [m]|692
Coverage [% of thickness]|97
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
