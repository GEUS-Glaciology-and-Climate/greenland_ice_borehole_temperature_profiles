Name|dye_3
Alternate name|DYE-3
Data source|Gundestrup, N. S., Hansen, B. Lyle: Bore-Hole Survey at Dye 3, South Greenland , Journal of Glaciology 30(106), Cambridge University Press (CUP), 282–288, 1984 
Drill year(s)|1979 to 1981
Data year(s)|1983
Longitude [°E]|-43.816667
Latitude [°N]|65.183333
Approximate location name|South Greenland
Location source|See data source
Ice thickness [m]|2038
Ice thickness year|1983
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|152
Depth of bottom measurement [m]|2030
