Name|devon_00
Alternate name|Devon borehole
Data source|WIC Email
Drill year(s)|1998-04-15 to 1998-05-07
Data year(s)|2000-04-15
Longitude [°E]|-82.14
Latitude [°N]|75.34
Approximate location name|Devon Ice Cap
Location source|
Ice thickness [m]|300.55
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|13
Depth of bottom measurement [m]|218
