Borehole ID|FOXX1
Place Name|FOXX
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|Lüthi, Martin P., Ryser, Claudia, Andrews, Lauren C., Catania, Ginny A., Funk, Martin, Hawley, Robert L., Hoffman, Matthew J., Neumann, Thomas A.: Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming , The Cryosphere 9(1), 245–253, 2015 
Data DOI|
Science Reference|Lüthi, M., C. Ryser, L. Andrews et al. 2015. Heat sources within the Greenland Ice Sheet: dissipation, temperate paleo-firn and cryo-hydrologic warming. The Cryosphere. 9: 245-253. 
Science DOI|10.5194/tc-9-245-2015
Date|2011-2013
Longitude [°E]|-49.8803
Latitude [°N]|69.4464
Location source|Colgan, 2021
Depth of top measurement [m]|6.0
Depth of bottom measurement [m]|611
Ice thickness [m]|631
Coverage [% of thickness]|96
Ice thickness source|Martin Luthi
General_Note|
Temperature_note|Digitized from graphic
Thickness_note|
Location_note|
