Borehole ID|Bowdoin_BH1
Place name|Bowdoin Glacier
Geographic location|Northwest Greenland
Site type|Ice sheet
Data Source|Seguinot, Funk, Bauder, Wyder, Senn, & Sugiyama. (2020). Bowdoin Glacier borehole temperature data [Data set]. Zenodo. https://doi.org/10.5281/zenodo.3695961
Data DOI|10.5281/zenodo.3695961
Science Source|Seguinot J, Funk M, Bauder A, Wyder T, Senn C and Sugiyama S (2020) Englacial Warming Indicates Deep Crevassing in Bowdoin Glacier, Greenland. Front. Earth Sci. 8:65. doi: 10.3389/feart.2020.00065
Science DOI|10.3389/feart.2020.00065
Date|2014-10-01
Longitude [°E]|-68.5565598058807
Latitude [°N]|77.69072896854759
Location Source|https://github.com/juseg/bowdoin/commit/aef3510
Depth of top measurement [m]|123.0
Depth of bottom measurement [m]|265
Ice thickness [m]|272
Coverage [% of thickness]|52
Ice thickness source|10.3389/feart.2020.00065
Note|
