Name|gisp2
Alternate name|GISP2; GISP II
Data source|Joe MacGregor email
Drill year(s)|
Data year(s)|1989,1990
Longitude [°E]|
Latitude [°N]|
Approximate location name|
Location source|
Ice thickness [m]|3100
Ice thickness year|
Ice thickness source|Hodge 1990?
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|100
Depth of bottom measurement [m]|3048
