Borehole ID|TD2_88
Place name|Paakitsoq
Geographic location|Central West Greenland
Site type|Ice sheet
Data Source|Lüthi email
Data DOI|
Science Source|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1988-05-19
Longitude [°E]|-50.1
Latitude [°N]|69.45
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|27.0
Depth of bottom measurement [m]|202
Ice thickness [m]|470
Coverage [% of thickness]|37
Ice thickness source|Unknown PDF: See td1
Note|
