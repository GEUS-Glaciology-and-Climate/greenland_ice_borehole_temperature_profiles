Name|grip
Alternate name|GRIP
Data source|Gary Clow email
Drill year(s)|1989-1992 (Vinther, 2008)
Data year(s)|
Longitude [°E]|-37.64
Latitude [°N]|72.58
Approximate location name|
Location source|Vinther (2008)
Ice thickness [m]|3028.57
Ice thickness year|
Ice thickness source|Data from Gary Clow
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|40.93
Depth of bottom measurement [m]|3028.57
