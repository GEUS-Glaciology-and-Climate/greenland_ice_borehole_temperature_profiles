Name|m2020_15s
Alternate name|
Data source|McDowell, Ian E., Humphrey, Neil F., Harper, Joel T., Meierbachtol, Toby W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet , The Cryosphere Discussions (In Review) , Copernicus GmbH, 8 2020 
Drill year(s)|
Data year(s)|2017
Longitude [°E]|
Latitude [°N]|
Approximate location name|
Location source|
Ice thickness [m]|660
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|B
Depth of top measurement [m]|35.0
Depth of bottom measurement [m]|655.0
