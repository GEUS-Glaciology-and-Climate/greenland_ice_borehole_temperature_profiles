Borehole ID|td3
Descriptive Name|
Area|Paakitsoq
Data reference|Unknown PDF: See td1. Also Phillips (2010)
Data DOI|
Science reference|
Science DOI|
Date|1988-08-18
Longitude [°E]|-50.0
Latitude [°N]|69.483
Location source|Unknown PDF: See td1. Also Phillips (2010)
Depth of top measurement [m]|20.0
Depth of bottom measurement [m]|350.0
Ice thickness [m]|350
Coverage [% of thickness]|94
Ice thickness source|Unknown PDF: See td1. Also Phillips (2010)
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
