Name|agassiz77
Alternate name|Agassiz 77 borehole 
Data source|WIC Email
Data year(s)|1977
Depth of top measurement [m]|11.0 
Depth of bottom measurement [m]|341.0 
Drill year(s)|1977 (Vinther, 2008)
Longitude [°E]|-73.1 
Latitude [°N]|80.7 
Approximate location name|Agassiz Ice Cap 
Location source|Vinther, 2008
Ice thickness [m]|340.9 
Ice thickness year|
Ice thickness source|See data source 
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|T 
