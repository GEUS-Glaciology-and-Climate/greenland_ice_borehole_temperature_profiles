Borehole ID|Agassiz84
Place Name|Agassiz Ice Cap
Geographic Location|Canadian Arctic North
Ice Type|Ice cap
Data Reference|W. Colgan email
Data DOI|
Science Reference|Clarke, G. K. C., Fisher, D. A., Waddington, E. D.: Wind pumping: A potentially significant heat source in ice sheets , The Physical Basis of Ice Sheet Modelling in Proceedings of the Vancouver Symposium, IAHS , volume 170, 169–180, 1987
Science DOI|
Date|1984
Longitude [°E]|-73.1
Latitude [°N]|80.7
Location source|Vinther, 2008
Depth of top measurement [m]|3.0
Depth of bottom measurement [m]|128
Ice thickness [m]|128
Coverage [% of thickness]|98
Ice thickness source|See data source
General_Note|
Temperature_note|
Thickness_note|Ice thickness from data does not match ice thickness from Vinther (2008)
Location_note|Location approximate
