Borehole ID|Store_S30
Place name|Store Glacier
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Doyle, S., B. Hubbard, P. Christoffersen, T. Young, C. Hofstede, M. Bougamont et al. (2018): SAFIRE borehole, AWS and GPS datasets. 
Data DOI|10.6084/m9.figshare.5745294.v1
Science Source|Doyle, S.H., Hubbard, B., Christoffersen, P., Young, T. J., Hofstede, C., Bougamont, M., Box, J. E. & Hubbard, A. 2018. Physical conditions of fast glacier flow: 1. Measurements from boreholes drilled to the bed of Store Glacier, West Greenland, Journal of Geophysical Research: Earth Surface, DOI: 10.1002/2017JF004529.
Science DOI|10.1002/2017JF004529
Date|2014
Longitude [°E]|-49.9167
Latitude [°N]|70.5167
Location Source|Doyle, 2018
Depth of top measurement [m]|102.0
Depth of bottom measurement [m]|604
Ice thickness [m]|600
Coverage [% of thickness]|84
Ice thickness source|Doyle (2018)
Velocity [m/yr]|598.3
Note|
