Name|mcdowell_2021_14w
Alternate name|
Data source| McDowell, I. E., Humphrey, N. F., Harper, J. T., and Meierbachtol, T. W.: The cooling signature of basal crevasses in a hard-bedded region of the Greenland Ice Sheet, The Cryosphere, 15, 897–907, https://doi.org/10.5194/tc-15-897-2021, 2021.
Drill year(s)|2014
Data year(s)|August 2015
Longitude [°E]|-49.57478802
Latitude [°N]|67.18201398
Approximate location name|
Location source|
Ice thickness [m]|661
Ice thickness year|2014
Ice thickness source|See raw data file `Greenland_AblationZone_TProfiles.xlsx` in 14n folder
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|B
Depth of top measurement [m]|40
Depth of bottom measurement [m]|660
