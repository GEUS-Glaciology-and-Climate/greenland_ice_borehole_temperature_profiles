Borehole ID|penny
Descriptive Name|Penny Ice Cap
Area|
Data reference|W. Colgan email
Data DOI|
Science reference|
Science DOI|
Date|1996
Longitude [°E]|-65.2
Latitude [°N]|67.3
Location source|
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|176.0
Ice thickness [m]|176
Coverage [% of thickness]|94
Ice thickness source|Data file + WIC email (see also Fisher 1998)
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
