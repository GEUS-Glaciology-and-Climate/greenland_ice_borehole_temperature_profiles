Borehole ID|TD2_88
Place Name|Paakitsoq
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|Unknown PDF: See td1
Data DOI|
Science Reference|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1988-05-19
Longitude [°E]|-50.1
Latitude [°N]|69.45
Location source|Colgan, 2021
Depth of top measurement [m]|27.0
Depth of bottom measurement [m]|202.0
Ice thickness [m]|470
Coverage [% of thickness]|37
Ice thickness source|Unknown PDF: See td1
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
