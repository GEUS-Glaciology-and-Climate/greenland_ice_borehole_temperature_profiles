Name|agassiz84
Alternate name|Agassiz 1984 borehole
Data source|WIC Email
Drill year(s)|nan
Data year(s)|1984
Longitude [°E]|-73.1
Latitude [°N]|80.7
Approximate location name|Agassiz Ice Cap
Location source|See data source
Ice thickness [m]|127.6
Ice thickness year|nan
Ice thickness source|See data source
Surface velocity [m yr^-1]|nan
Surface velocity year|nan
Surface velocity source|nan
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|3.0
Depth of bottom measurement [m]|128.0
Coverage [% of thickness]|98
