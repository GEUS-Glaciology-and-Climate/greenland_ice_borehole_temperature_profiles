Borehole ID|Isunnguata_13km-10
Place name|Isunnguata Sermia
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Meierbachtol email
Data DOI|
Science Source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A941
Date|2010
Longitude [°E]|-50.02945
Latitude [°N]|67.19158
Location Source|T. Meierbachtol email
Depth of top measurement [m]|4.0
Depth of bottom measurement [m]|559
Ice thickness [m]|704
Coverage [% of thickness]|79
Ice thickness source|BedMachine v4
Note|See data in M1-10 folder; Harrington 2015 name: S2
