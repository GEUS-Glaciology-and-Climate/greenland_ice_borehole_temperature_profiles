Borehole ID|Store_R29
Place name|Store Glacier
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Hubbard, Bryn; Christoffersen, Poul; Doyle, Samuel; Chudley, Thomas; Schoonman, Charlotte; Law, Robert; et al. (2020): Supporting data for 'Borehole-based characterization of deep crevasses at a Greenlandic outlet glacier' published in AGU Advances. figshare. Dataset. https://doi.org/10.6084/m9.figshare.13400072.v1
Data DOI|10.6084/m9.figshare.13400072.v2
Science Source|Hubbard, B., Christoffersen, P., Doyle, S. H., Chudley, T. R., Bougamont, M. H., Law, R., & Schoonman, C. (2020). Borehole-based characterization of deep crevasses at a Greenlandic outlet glacier.
Science DOI|10.1029/2020AV000291
Date|2018-08
Longitude [°E]|-50.05894
Latitude [°N]|70.56359
Location Source|S. Doyle email
Depth of top measurement [m]|27.0
Depth of bottom measurement [m]|949
Ice thickness [m]|949
Coverage [% of thickness]|97
Ice thickness source|See science reference
Note|Note: Temperature measured in immediately adjacent Boreholes 18b and 18d.
