Borehole ID|GULL
Place name|Sermeq Avannerleq
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Ryser, C., Lüthi, M. P., Andrews, L. C., Hoffman, M. J., Catania, G. A., Hawley, R. L., ... & Kristensen, S. S. (2014). Sustained high basal motion of the Greenland ice sheet revealed by borehole deformation. Journal of Glaciology, 60(222), 647-660.
Data DOI|10.3189/2014JoG13J196
Science Source|Ryser, C., Lüthi, M. P., Andrews, L. C., Hoffman, M. J., Catania, G. A., Hawley, R. L., ... & Kristensen, S. S. (2014). Sustained high basal motion of the Greenland ice sheet revealed by borehole deformation. Journal of Glaciology, 60(222), 647-660.
Science DOI|10.3189/2014JoG13J196
Date|2012
Longitude [°E]|-49.7182
Latitude [°N]|69.4524
Location Source|10.3189/2014JoG13J196
Depth of top measurement [m]|4.0
Depth of bottom measurement [m]|705
Ice thickness [m]|705
Coverage [% of thickness]|99
Ice thickness source|Ryser, 2014 (Table 3). 705/707 for thickness
Note|Only using 'string1' near bottom. Date: Data was collected in 2011 and 2012 and the data extracted from the cooling curves
