Name|agassiz79b
Alternate name|Agassiz ice cap 1979B borehole
Data source|WIC Email
Drill year(s)|1979 (Vinther, 2008)
Data year(s)|1979
Longitude [°E]|-73.1
Latitude [°N]|80.7
Approximate location name|Agassiz Ice Cap
Location source|Vinther (2008)
Ice thickness [m]|141.2
Ice thickness year|nan
Ice thickness source|See data source
Surface velocity [m yr^-1]|nan
Surface velocity year|nan
Surface velocity source|nan
Measured from: Top, Bottom, Relative|T
Depth of top measurement [m]|11.0
Depth of bottom measurement [m]|141.0
Coverage [% of thickness]|92
