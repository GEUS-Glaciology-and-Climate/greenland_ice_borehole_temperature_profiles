Name|tuto_ramp
Alternate name|Tuto Ramp
Data source|Davis, RM: Approach roads, Greenland 1960–1964 , Technical Report 133. Corps of Engineers, Cold Regions Research & Engineering Laboratory , 1967 
Data year(s)|1962 (August)
Depth of top measurement [m]|
Depth of bottom measurement [m]|
Drill year(s)|
Longitude [°E]|-68.287295
Latitude [°N]|76.41133
Approximate location name|Thule Approach Road(?)
Location source|
Ice thickness [m]|48
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|1.0
Surface velocity year|
Surface velocity source|WIC Email
Measured from: Top, Bottom, Relative|T(ish)
