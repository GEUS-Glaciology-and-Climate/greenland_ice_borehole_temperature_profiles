Name|hanstausen_hare
Alternate name|Hans Tausen Hare
Data source|Zekollari, Harry, Huybrechts, Philippe, Noël, Brice, van de Berg, Willem Jan, van den Broeke, Michiel R.: Sensitivity, stability and future evolution of the world’s northernmost ice cap, Hans Tausen Iskappe (Greenland) , The Cryosphere 11(2), Copernicus GmbH, 805–825, 3 2017 
Drill year(s)|
Data year(s)|
Longitude [°E]|
Latitude [°N]|
Approximate location name|
Location source|
Ice thickness [m]|289
Ice thickness year|
Ice thickness source|See data source
Surface velocity [m yr^-1]|
Surface velocity year|
Surface velocity source|
Measured from: Top, Bottom, Relative|B
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|288.0
