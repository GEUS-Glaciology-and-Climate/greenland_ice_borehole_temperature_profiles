Borehole ID|Jakobshavn95D_T4
Place Name|Jakobshavn Isbræ
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|M. Lüthi email
Data DOI|
Science Reference|Lüthi, Martin, Funk, Martin, Iken, Almut, Gogineni, Shivaprasad, Truffer, Martin: Mechanisms of fast flow in Jakobshavns Isbræ, West Greenland: Part III. Measurements of ice deformation, temperature and cross-borehole conductivity in boreholes to the bedrock, Journal of Glaciology 48(162), 369–385, 2002 
Science DOI|10.3189/172756502781831322
Date|1995
Longitude [°E]|-48.6871
Latitude [°N]|69.235
Location source|Colgan, 2021
Depth of top measurement [m]|450.0
Depth of bottom measurement [m]|600.0
Ice thickness [m]|832
Coverage [% of thickness]|18
Ice thickness source|See science reference
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|Location from Geothermal Database
