Borehole ID|StationCentrale
Place Name|Station Centrale
Geographic Location|Northwest Greenland
Ice Type|Ice sheet
Data Reference|Heuberger, J.-C. 1954. Expéditions Polaires Françaises: Missions Paul-Emil Victor. Glaciologie Groenland Volume 1: Forages sur l'inlandsis. Hermann & Cle, Éditeurs. Paris.
Data DOI|
Science Reference|Heuberger, J.-C. 1954. Expéditions Polaires Françaises: Missions Paul-Emil Victor. Glaciologie Groenland Volume 1: Forages sur l'inlandsis. Hermann & Cle, Éditeurs. Paris.
Science DOI|
Date|
Longitude [°E]|
Latitude [°N]|
Location source|
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|150
Ice thickness [m]|
Coverage [% of thickness]|#DIV/0!
Ice thickness source|
General_Note|
Temperature_note|https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/files/7082104/heuberger_1954.pdf
Thickness_note|
Location_note|
