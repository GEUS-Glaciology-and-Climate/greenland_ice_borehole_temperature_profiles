Borehole ID|td41
Descriptive Name|
Area|Paakitsoq
Data reference|Unknown PDF: See td1
Data DOI|
Science reference|
Science DOI|
Date|1991-11-05
Longitude [°E]|-49.683
Latitude [°N]|69.533
Location source|Unknown PDF: See td1
Depth of top measurement [m]|5.0
Depth of bottom measurement [m]|495.0
Ice thickness [m]|>600
Coverage [% of thickness]|#VALUE!
Ice thickness source|Unknown PDF: See td1
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
