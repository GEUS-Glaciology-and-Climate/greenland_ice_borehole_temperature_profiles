Borehole ID|Isua_11
Place name|Isua
Geographic location|Central West Greenland
Site type|Ice sheet
Data Source|Graphic in science source
Data DOI|
Science Source|Colebeck, S. and A. Gow. 1979. The margin of the Greenland Ice Sheet at Isua. Journal of Glaciology. 24: 155-165. 
Science DOI|10.3189/S0022143000014714
Date|1973
Longitude [°E]|-49.751
Latitude [°N]|65.2072
Location Source|10.5194/essd-2021-290
Depth of top measurement [m]|25.0
Depth of bottom measurement [m]|116
Ice thickness [m]|120
Coverage [% of thickness]|76
Ice thickness source|See data source
Note|"Measuremnet date 1972 or 1973. From Colbeck (1979), ""Five holes (see Fig. 3) were drilled in 1972 and 1973 for the purpose of making temperature measurements and taking ice cores."""
