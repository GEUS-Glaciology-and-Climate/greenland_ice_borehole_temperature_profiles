Borehole ID|pow
Descriptive Name|Prince of Wales
Area|
Data reference|W. Colgan email
Data DOI|
Science reference|
Science DOI|
Date|2005-05-15
Longitude [°E]|-80.395
Latitude [°N]|78.3897
Location source|
Depth of top measurement [m]|10.0
Depth of bottom measurement [m]|176.0
Ice thickness [m]|176
Coverage [% of thickness]|94
Ice thickness source|WIC
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
