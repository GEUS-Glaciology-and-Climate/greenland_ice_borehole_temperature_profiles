Borehole ID|TD4_91a
Place Name|Paakitsoq
Geographic Location|Central West Greenland
Ice Type|Ice sheet
Data Reference|Unknown PDF: See td1
Data DOI|
Science Reference|Thomsen, H.H., O.B. Olesen, R.J. Braithwaite, and C.E. Bøggild. 1991. Ice drilling and mass balance at Pakitsoq, Jakobshavn, central West Greenland. Rapport Grønlands Geologiske Undersøgelse, 152, 80–84. 
Science DOI|10.34194/rapggu.v152.8160
Date|1991-11-05
Longitude [°E]|-49.68
Latitude [°N]|69.53
Location source|Colgan, 2021
Depth of top measurement [m]|5.0
Depth of bottom measurement [m]|495
Ice thickness [m]|660
Coverage [% of thickness]|74
Ice thickness source|Estimate from Martin Luthi
General_Note|
Temperature_note|See https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/blob/main/TD1_88/Shallow88II.pdf and https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/blob/main/TD1_88/Thomsen_TD1_TD2_TD3_records.pdf
Thickness_note|
Location_note|
