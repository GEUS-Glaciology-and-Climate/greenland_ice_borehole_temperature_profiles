Borehole ID|Isunnguata_46km-11B
Place Name|Isunnguata Sermia
Geographic Location|Central West Greenland
Ice Type|
Data Reference|T. Meierbachtol email
Data DOI|
Science Reference|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A949
Date|2011
Longitude [°E]|-49.2891
Latitude [°N]|67.20134
Location source|T. Meierbachtol email
Depth of top measurement [m]|114.0
Depth of bottom measurement [m]|728.0
Ice thickness [m]|815.0
Coverage [% of thickness]|75
Ice thickness source|T. Meierbachtol email
Measured from: Top, Bottom, Relative|T
General_Note|See data in M1-10 folder
Temperature_note|
Thickness_note|
Location_note|Harrington 2015 name: S5-B
