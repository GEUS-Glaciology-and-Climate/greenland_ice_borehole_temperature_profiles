Borehole ID|Isunnguata_27km-11B
Place name|Isunnguata Sermia
Geographic location|Central West Greenland
Ice type|Ice sheet
Data Source|Meierbachtol email
Data DOI|
Science Source|Harrington, Joel A., Humphrey, Neil F., Harper, Joel T.: Temperature distribution and thermal anomalies along a flowline of the Greenland ice sheet , Annals of Glaciology 56(70), 98–104, 2015 
Science DOI|10.3189/2015AoG70A943
Date|2011
Longitude [°E]|-49.71913
Latitude [°N]|67.19527
Location Source|Meierbachtol email
Depth of top measurement [m]|27.0
Depth of bottom measurement [m]|460
Ice thickness [m]|466
Coverage [% of thickness]|93
Ice thickness source|T. Meierbachtol email
Velocity [m/yr]|98.7
Note|See data in M1-10 folder; Harrington 2015 name: S3-B
