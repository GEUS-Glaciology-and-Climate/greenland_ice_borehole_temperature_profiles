Borehole ID|SomeID
Place name|Some Glacier
Geographic location|Some Place
Site type|...
Data Source|An email or some reference
Data DOI|
Science Source|Reference
Science DOI|DOI
Date|YYYY-MM-DD
Longitude [°E]|-42.42
Latitude [°N]|42.42
Location Source|DOI
Depth of top measurement [m]|num
Depth of bottom measurement [m]|num
Ice thickness [m]|num
Coverage [% of thickness]|num
Ice thickness source|DOI or refenece or "See data source"
Note|Anything else
