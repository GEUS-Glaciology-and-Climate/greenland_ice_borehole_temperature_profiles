Borehole ID|StationCentrale_EGIG
Place Name|Station Centrale
Geographic Location|Northwest Greenland
Ice Type|Ice sheet
Data Reference|Brockamp, 1959
Data DOI|
Science Reference|
Science DOI|
Date|1959
Longitude [°E]|-56.07
Latitude [°N]|76.98
Location source|Colgan, 2021
Depth of top measurement [m]|20.0
Depth of bottom measurement [m]|150
Ice thickness [m]|
Coverage [% of thickness]|#DIV/0!
Ice thickness source|BedMachine_V3
General_Note|
Temperature_note|Digitized from https://github.com/GEUS-Glaciology-and-Climate/greenland_ice_borehole_temperature_profiles/files/7185520/Polarforsch1965_1-2_8.pdf
Thickness_note|Assuming same location as StationCentrale
Location_note|Assuming same location as StationCentrale
