Borehole ID|Isua_13
Place Name|Isua
Geographic Location|Central West Greenland
Ice Type|
Data Reference|Colbeck, S. C., Gow, A. J.: The Margin of the Greenland Ice Sheet at Isua , Journal of Glaciology 24(90), Cambridge University Press (CUP), 155–165, 1979 
Data DOI|
Science Reference|Colebeck, S. and A. Gow. 1979. The margin of the Greenland Ice Sheet at Isua. Journal of Glaciology. 24: 155-165. 
Science DOI|10.3189/S0022143000014714
Date|1972-1973
Longitude [°E]|-49.7456
Latitude [°N]|65.2069
Location source|Colgan2021
Depth of top measurement [m]|6.0
Depth of bottom measurement [m]|247.0
Ice thickness [m]|265.0
Coverage [% of thickness]|91
Ice thickness source|See data source
Measured from: Top, Bottom, Relative|T
General_Note|
Temperature_note|
Thickness_note|
Location_note|
